library ieee;
use ieee.std_logic_1164.all;

library work;
use work.types.all;

package sprites is
type palette_ROM is array (0 to 127) of std_logic_vector(7 downto 0);

constant red_rom : palette_ROM := (
x"fa",x"d2",x"e9",x"9b",x"ff",x"e4",x"a4",x"cd",
x"94",x"b5",x"d6",x"df",x"d1",x"c3",x"75",x"6a",
x"e6",x"84",x"ab",x"e4",x"ba",x"54",x"a1",x"b5",
x"b1",x"c5",x"dc",x"68",x"f0",x"e1",x"d0",x"62",
x"52",x"5b",x"c8",x"d9",x"59",x"5b",x"d5",x"62",
x"dc",x"52",x"5d",x"f5",x"f7",x"69",x"5c",x"da",
x"e2",x"e3",x"f3",x"67",x"e9",x"d9",x"d6",x"ee",
x"55",x"5d",x"db",x"8d",x"b1",x"96",x"df",x"df",
x"d9",x"c9",x"c0",x"4e",x"d9",x"de",x"5a",x"60",
x"5d",x"de",x"8d",x"5e",x"5e",x"79",x"df",x"5a",
x"68",x"5e",x"c9",x"ff",x"ed",x"58",x"14",x"fc",
x"fc",x"73",x"9c",x"00",x"ec",x"fc",x"d3",x"f0",
x"fd",x"d7",x"00",x"ff",x"ed",x"e9",x"f9",x"5d",
x"c7",x"ff",x"d6",x"e4",x"d9",x"e3",x"9e",x"d0",
x"84",x"b9",x"87",x"f8",x"bd",x"ef",x"ea",x"4f",
x"e0",x"fc",x"fa",x"5d",x"ac",x"fc",x"d7",x"ff");

constant green_rom : palette_ROM := (
x"fa",x"ef",x"fc",x"da",x"28",x"e4",x"c6",x"ec",
x"b7",x"d4",x"d6",x"df",x"ec",x"e0",x"9c",x"ca",
x"fa",x"a9",x"e3",x"fd",x"e7",x"38",x"dc",x"e5",
x"e5",x"eb",x"ee",x"91",x"f0",x"f9",x"ed",x"cc",
x"c3",x"cb",x"c0",x"ed",x"de",x"e1",x"f0",x"df",
x"f6",x"cb",x"c7",x"f5",x"f7",x"cd",x"de",x"f7",
x"f1",x"fa",x"f3",x"df",x"e9",x"d9",x"f4",x"ee",
x"80",x"87",x"f6",x"d8",x"e4",x"d8",x"f0",x"f9",
x"f3",x"e5",x"dd",x"c0",x"f4",x"f8",x"84",x"8a",
x"88",x"d8",x"b1",x"e2",x"df",x"a0",x"f9",x"df",
x"90",x"df",x"e6",x"ff",x"ed",x"d8",x"18",x"fc",
x"a0",x"bf",x"e6",x"00",x"ec",x"78",x"ce",x"ea",
x"fd",x"a8",x"a8",x"b1",x"f2",x"e1",x"f7",x"e2",
x"c2",x"db",x"be",x"60",x"97",x"c3",x"98",x"ce",
x"7f",x"81",x"86",x"b7",x"a2",x"ed",x"a2",x"c1",
x"80",x"38",x"d7",x"e1",x"cc",x"e0",x"e6",x"ff");

constant blue_rom : palette_ROM := (
x"fa",x"c6",x"d9",x"d5",x"09",x"e4",x"5c",x"c4",
x"51",x"68",x"d6",x"df",x"7d",x"73",x"3a",x"cd",
x"d8",x"45",x"ba",x"8b",x"c3",x"47",x"d7",x"c4",
x"bc",x"bc",x"cf",x"30",x"f0",x"d8",x"c8",x"7c",
x"cb",x"78",x"c0",x"cf",x"6e",x"6f",x"c6",x"76",
x"85",x"6c",x"cc",x"f5",x"f7",x"7f",x"71",x"d8",
x"d0",x"d8",x"f3",x"77",x"e9",x"d9",x"d7",x"ee",
x"22",x"28",x"85",x"c9",x"c5",x"cf",x"cf",x"87",
x"83",x"77",x"71",x"ca",x"83",x"d8",x"26",x"2a",
x"28",x"95",x"4b",x"70",x"70",x"3d",x"88",x"6f",
x"2f",x"72",x"78",x"ff",x"ed",x"58",x"1c",x"fc",
x"48",x"2e",x"59",x"00",x"ec",x"58",x"8e",x"a1",
x"fd",x"4c",x"48",x"41",x"61",x"e1",x"f7",x"70",
x"86",x"5f",x"9b",x"18",x"37",x"55",x"98",x"ce",
x"7f",x"2f",x"86",x"33",x"47",x"ed",x"3c",x"ca",
x"2c",x"00",x"8c",x"6f",x"62",x"b4",x"cc",x"ff");

type flappy_rom is array (0 to 2, 0 to BirdWidth, 0 to BirdHeight) of integer range 0 to 127;
constant flappy_bird : flappy_rom := ((
(127,127,127,127,127,127,127,127,21,21,21,21,21,21,127,127,127,127,127,127,127,127,127,127),
(127,127,127,127,127,127,127,127,21,21,21,21,21,21,127,127,127,127,127,127,127,127,127,127),
(127,127,127,127,127,127,21,21,0,0,0,0,122,122,21,21,127,127,127,127,127,127,127,127),
(127,127,127,127,127,127,21,21,0,0,0,0,122,122,21,21,127,127,127,127,127,127,127,127),
(127,127,127,127,127,127,21,21,0,0,0,0,0,0,122,122,21,21,21,21,127,127,127,127),
(127,127,127,127,127,127,21,21,0,0,0,0,0,0,122,122,21,21,21,21,127,127,127,127),
(127,127,127,127,21,21,21,21,0,0,0,0,0,0,122,122,21,21,120,120,21,21,127,127),
(127,127,127,127,21,21,21,21,0,0,0,0,0,0,122,122,21,21,120,120,21,21,127,127),
(127,127,21,21,122,122,21,21,0,0,0,0,0,0,122,122,21,21,120,120,21,21,127,127),
(127,127,21,21,122,122,21,21,0,0,0,0,0,0,122,122,21,21,120,120,21,21,127,127),
(127,127,21,21,122,122,115,115,21,21,0,0,122,122,21,21,120,120,120,120,120,120,21,21),
(127,127,21,21,122,122,115,115,21,21,0,0,122,122,21,21,120,120,120,120,120,120,21,21),
(21,21,122,122,115,115,115,115,115,115,21,21,21,21,115,115,120,120,120,120,120,120,21,21),
(21,21,122,122,115,115,115,115,115,115,21,21,21,21,115,115,120,120,120,120,120,120,21,21),
(21,21,122,122,115,115,115,115,115,115,115,115,115,115,115,115,120,120,120,120,120,120,21,21),
(21,21,122,122,115,115,115,115,115,115,115,115,115,115,115,115,120,120,120,120,120,120,21,21),
(21,21,122,122,21,21,21,21,21,21,115,115,115,115,115,115,21,21,120,120,120,120,21,21),
(21,21,122,122,21,21,21,21,21,21,115,115,115,115,115,115,21,21,120,120,120,120,21,21),
(21,21,21,21,0,0,126,126,126,126,21,21,115,115,21,21,121,121,21,21,120,120,21,21),
(21,21,21,21,0,0,126,126,126,126,21,21,115,115,21,21,121,121,21,21,120,120,21,21),
(21,21,0,0,0,0,0,0,0,0,126,126,21,21,121,121,21,21,121,121,21,21,127,127),
(21,21,0,0,0,0,0,0,0,0,126,126,21,21,121,121,21,21,121,121,21,21,127,127),
(21,21,0,0,0,0,0,0,0,0,0,0,21,21,121,121,21,21,121,121,21,21,127,127),
(21,21,0,0,0,0,0,0,0,0,0,0,21,21,121,121,21,21,121,121,21,21,127,127),
(127,127,21,21,0,0,21,21,21,21,0,0,21,21,121,121,21,21,121,121,21,21,127,127),
(127,127,21,21,0,0,21,21,21,21,0,0,21,21,121,121,21,21,121,121,21,21,127,127),
(127,127,127,127,21,21,0,0,0,0,0,0,21,21,121,121,21,21,121,121,21,21,127,127),
(127,127,127,127,21,21,0,0,0,0,0,0,21,21,121,121,21,21,121,121,21,21,127,127),
(127,127,127,127,127,127,21,21,21,21,21,21,21,21,121,121,21,21,121,121,21,21,127,127),
(127,127,127,127,127,127,21,21,21,21,21,21,21,21,121,121,21,21,121,121,21,21,127,127),
(127,127,127,127,127,127,127,127,127,127,127,127,21,21,121,121,21,21,21,21,127,127,127,127),
(127,127,127,127,127,127,127,127,127,127,127,127,21,21,121,121,21,21,21,21,127,127,127,127),
(127,127,127,127,127,127,127,127,127,127,127,127,127,127,21,21,127,127,127,127,127,127,127,127),
(127,127,127,127,127,127,127,127,127,127,127,127,127,127,21,21,127,127,127,127,127,127,127,127)
),(
(127,127,127,127,127,127,127,127,127,127,127,127,21,21,21,21,127,127,127,127,127,127,127,127),
(127,127,127,127,127,127,127,127,127,127,127,127,21,21,21,21,127,127,127,127,127,127,127,127),
(127,127,127,127,127,127,127,127,21,21,21,21,0,0,122,122,21,21,127,127,127,127,127,127),
(127,127,127,127,127,127,127,127,21,21,21,21,0,0,122,122,21,21,127,127,127,127,127,127),
(127,127,127,127,127,127,21,21,115,115,21,21,0,0,0,0,21,21,21,21,127,127,127,127),
(127,127,127,127,127,127,21,21,115,115,21,21,0,0,0,0,21,21,21,21,127,127,127,127),
(127,127,127,127,21,21,122,122,115,115,21,21,0,0,0,0,21,21,120,120,21,21,127,127),
(127,127,127,127,21,21,122,122,115,115,21,21,0,0,0,0,21,21,120,120,21,21,127,127),
(127,127,21,21,122,122,115,115,115,115,21,21,0,0,0,0,21,21,120,120,21,21,127,127),
(127,127,21,21,122,122,115,115,115,115,21,21,0,0,0,0,21,21,120,120,21,21,127,127),
(127,127,21,21,122,122,115,115,115,115,21,21,0,0,122,122,21,21,120,120,120,120,21,21),
(127,127,21,21,122,122,115,115,115,115,21,21,0,0,122,122,21,21,120,120,120,120,21,21),
(21,21,122,122,115,115,115,115,115,115,115,115,21,21,21,21,120,120,120,120,120,120,21,21),
(21,21,122,122,115,115,115,115,115,115,115,115,21,21,21,21,120,120,120,120,120,120,21,21),
(21,21,122,122,115,115,115,115,115,115,115,115,115,115,115,115,120,120,120,120,120,120,21,21),
(21,21,122,122,115,115,115,115,115,115,115,115,115,115,115,115,120,120,120,120,120,120,21,21),
(21,21,122,122,21,21,21,21,21,21,115,115,115,115,115,115,21,21,120,120,120,120,21,21),
(21,21,122,122,21,21,21,21,21,21,115,115,115,115,115,115,21,21,120,120,120,120,21,21),
(21,21,21,21,0,0,126,126,126,126,21,21,115,115,21,21,121,121,21,21,120,120,21,21),
(21,21,21,21,0,0,126,126,126,126,21,21,115,115,21,21,121,121,21,21,120,120,21,21),
(21,21,0,0,0,0,0,0,0,0,126,126,21,21,121,121,21,21,121,121,21,21,127,127),
(21,21,0,0,0,0,0,0,0,0,126,126,21,21,121,121,21,21,121,121,21,21,127,127),
(21,21,0,0,0,0,0,0,0,0,0,0,21,21,121,121,21,21,121,121,21,21,127,127),
(21,21,0,0,0,0,0,0,0,0,0,0,21,21,121,121,21,21,121,121,21,21,127,127),
(127,127,21,21,0,0,21,21,21,21,0,0,21,21,121,121,21,21,121,121,21,21,127,127),
(127,127,21,21,0,0,21,21,21,21,0,0,21,21,121,121,21,21,121,121,21,21,127,127),
(127,127,127,127,21,21,0,0,0,0,0,0,21,21,121,121,21,21,121,121,21,21,127,127),
(127,127,127,127,21,21,0,0,0,0,0,0,21,21,121,121,21,21,121,121,21,21,127,127),
(127,127,127,127,127,127,21,21,21,21,21,21,21,21,121,121,21,21,121,121,21,21,127,127),
(127,127,127,127,127,127,21,21,21,21,21,21,21,21,121,121,21,21,121,121,21,21,127,127),
(127,127,127,127,127,127,127,127,127,127,127,127,21,21,121,121,21,21,21,21,127,127,127,127),
(127,127,127,127,127,127,127,127,127,127,127,127,21,21,121,121,21,21,21,21,127,127,127,127),
(127,127,127,127,127,127,127,127,127,127,127,127,127,127,21,21,127,127,127,127,127,127,127,127),
(127,127,127,127,127,127,127,127,127,127,127,127,127,127,21,21,127,127,127,127,127,127,127,127)),(
(127,127,127,127,127,127,127,127,127,127,127,127,127,127,21,21,21,21,21,21,127,127,127,127),
(127,127,127,127,127,127,127,127,127,127,127,127,127,127,21,21,21,21,21,21,127,127,127,127),
(127,127,127,127,127,127,127,127,21,21,21,21,21,21,122,122,0,0,0,0,21,21,127,127),
(127,127,127,127,127,127,127,127,21,21,21,21,21,21,122,122,0,0,0,0,21,21,127,127),
(127,127,127,127,127,127,21,21,115,115,115,115,21,21,0,0,0,0,0,0,21,21,127,127),
(127,127,127,127,127,127,21,21,115,115,115,115,21,21,0,0,0,0,0,0,21,21,127,127),
(127,127,127,127,21,21,122,122,115,115,115,115,21,21,0,0,0,0,122,122,21,21,127,127),
(127,127,127,127,21,21,122,122,115,115,115,115,21,21,0,0,0,0,122,122,21,21,127,127),
(127,127,21,21,122,122,115,115,115,115,115,115,21,21,0,0,0,0,21,21,21,21,127,127),
(127,127,21,21,122,122,115,115,115,115,115,115,21,21,0,0,0,0,21,21,21,21,127,127),
(127,127,21,21,122,122,115,115,115,115,115,115,21,21,122,122,21,21,120,120,120,120,21,21),
(127,127,21,21,122,122,115,115,115,115,115,115,21,21,122,122,21,21,120,120,120,120,21,21),
(21,21,122,122,115,115,115,115,115,115,115,115,115,115,21,21,120,120,120,120,120,120,21,21),
(21,21,122,122,115,115,115,115,115,115,115,115,115,115,21,21,120,120,120,120,120,120,21,21),
(21,21,122,122,115,115,115,115,115,115,115,115,115,115,115,115,120,120,120,120,120,120,21,21),
(21,21,122,122,115,115,115,115,115,115,115,115,115,115,115,115,120,120,120,120,120,120,21,21),
(21,21,122,122,21,21,21,21,21,21,115,115,115,115,115,115,21,21,120,120,120,120,21,21),
(21,21,122,122,21,21,21,21,21,21,115,115,115,115,115,115,21,21,120,120,120,120,21,21),
(21,21,21,21,0,0,126,126,126,126,21,21,115,115,21,21,121,121,21,21,120,120,21,21),
(21,21,21,21,0,0,126,126,126,126,21,21,115,115,21,21,121,121,21,21,120,120,21,21),
(21,21,0,0,0,0,0,0,0,0,126,126,21,21,121,121,21,21,121,121,21,21,127,127),
(21,21,0,0,0,0,0,0,0,0,126,126,21,21,121,121,21,21,121,121,21,21,127,127),
(21,21,0,0,0,0,0,0,0,0,0,0,21,21,121,121,21,21,121,121,21,21,127,127),
(21,21,0,0,0,0,0,0,0,0,0,0,21,21,121,121,21,21,121,121,21,21,127,127),
(127,127,21,21,0,0,21,21,21,21,0,0,21,21,121,121,21,21,121,121,21,21,127,127),
(127,127,21,21,0,0,21,21,21,21,0,0,21,21,121,121,21,21,121,121,21,21,127,127),
(127,127,127,127,21,21,0,0,0,0,0,0,21,21,121,121,21,21,121,121,21,21,127,127),
(127,127,127,127,21,21,0,0,0,0,0,0,21,21,121,121,21,21,121,121,21,21,127,127),
(127,127,127,127,127,127,21,21,21,21,21,21,21,21,121,121,21,21,121,121,21,21,127,127),
(127,127,127,127,127,127,21,21,21,21,21,21,21,21,121,121,21,21,121,121,21,21,127,127),
(127,127,127,127,127,127,127,127,127,127,127,127,21,21,121,121,21,21,21,21,127,127,127,127),
(127,127,127,127,127,127,127,127,127,127,127,127,21,21,121,121,21,21,21,21,127,127,127,127),
(127,127,127,127,127,127,127,127,127,127,127,127,127,127,21,21,127,127,127,127,127,127,127,127),
(127,127,127,127,127,127,127,127,127,127,127,127,127,127,21,21,127,127,127,127,127,127,127,127))
);

type bg_rom is array (0 to 287, 0 to 83) of integer range 0 to 127;
constant bg_bird : bg_rom := (
(67,67,67,67,67,67,67,67,67,119,119,42,42,15,15,29,29,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,29,29,22,22,60,60,3,3,60,23,20,23,20,20,23,20,20,20,20,20,23,23,23,23,3,3,61,61,59,59,31,33,39,39,37,37,75,75,75,75,75,75,75,75,75),
(67,67,67,67,67,67,67,67,67,119,119,32,42,15,15,29,29,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,29,29,22,3,60,60,3,3,23,23,23,20,20,20,20,20,20,20,20,20,20,20,23,23,3,3,61,61,59,59,33,33,39,39,37,37,75,75,75,75,75,75,75,75,75),
(67,67,67,67,67,67,67,119,119,32,32,15,15,47,47,49,49,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,29,29,22,22,30,30,3,3,30,30,1,1,1,1,1,1,1,1,1,1,1,1,1,1,30,30,7,7,25,25,31,31,39,39,123,123,75,75,75,75,75,75,75,75,75),
(67,67,67,67,67,67,67,119,119,32,32,15,42,47,47,49,49,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,29,29,22,22,7,30,3,3,30,30,1,1,38,1,1,1,1,1,1,1,1,1,1,1,30,30,7,7,25,25,31,31,39,39,123,123,75,75,75,75,75,75,75,75,75),
(67,67,67,67,67,67,67,32,32,42,42,54,54,29,29,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,49,49,22,22,22,3,3,3,30,1,1,1,20,20,20,20,38,38,20,20,20,20,1,1,22,22,3,3,25,25,45,45,51,51,123,123,103,103,103,103,103,103,103,103,75),
(67,67,67,67,67,67,67,32,32,42,42,54,54,29,29,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,49,49,22,22,22,22,22,22,30,1,1,1,20,20,20,20,38,38,20,20,20,20,1,1,22,22,3,22,25,7,31,45,51,51,123,123,103,103,103,103,103,103,103,103,75),
(67,67,67,67,67,119,119,32,32,15,15,69,47,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,29,49,69,69,22,22,1,1,38,38,38,38,38,38,38,38,38,38,38,38,38,38,1,1,7,7,25,25,25,25,41,33,76,76,37,37,37,37,37,37,123,123,103),
(67,67,67,67,67,119,119,32,32,15,15,47,69,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,29,29,69,69,22,22,1,1,38,38,38,38,38,38,38,38,38,38,38,38,38,38,1,1,1,7,25,7,25,25,33,33,76,76,37,37,37,37,37,37,123,123,103),
(67,67,67,67,67,32,32,42,42,54,54,29,29,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,29,29,22,22,1,1,1,1,20,20,20,20,1,1,20,20,20,20,1,1,3,22,61,3,25,25,31,33,41,41,79,46,79,79,79,79,41,41,37,37,103),
(67,67,67,67,67,32,32,42,42,54,54,29,29,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,29,29,22,22,1,1,1,1,20,20,20,20,1,1,20,20,20,20,1,1,22,3,3,3,25,25,31,31,41,33,36,46,79,79,79,79,41,41,37,37,103),
(67,67,67,119,119,32,32,15,15,69,47,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,29,29,22,22,30,30,30,30,1,1,1,1,1,1,1,1,1,1,30,30,7,7,25,25,45,45,51,51,81,46,41,41,36,36,41,41,79,37,37,37,103),
(67,67,67,119,119,32,32,15,15,47,69,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,29,29,22,22,38,1,30,30,38,1,1,1,1,1,1,1,1,1,30,30,7,7,25,25,45,45,51,51,46,81,41,41,36,36,41,41,79,79,37,37,103),
(67,67,67,119,119,42,42,54,54,29,29,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,49,49,22,22,22,22,22,22,22,22,22,22,22,22,22,22,22,22,22,22,3,61,59,59,33,33,81,39,79,79,41,41,36,36,41,41,37,37,123,123,75),
(67,67,67,119,119,42,32,54,54,29,29,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,49,49,22,22,22,22,22,22,22,22,22,22,22,22,22,22,22,22,3,22,61,3,59,59,33,33,39,81,79,79,41,41,36,36,41,41,37,37,123,123,75),
(67,67,67,32,32,42,42,47,47,49,49,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,49,16,26,62,26,26,26,26,26,26,26,26,26,26,26,26,35,35,7,30,45,45,39,51,81,46,37,37,79,79,41,41,79,79,37,37,103,103,75),
(67,67,67,32,32,42,42,47,54,49,49,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,49,49,26,26,26,26,26,26,26,26,26,26,26,26,26,26,35,35,7,7,31,45,39,39,81,103,37,37,79,79,41,41,79,79,37,37,103,103,75),
(67,67,67,32,32,42,42,69,47,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,62,48,62,62,62,62,62,62,62,62,62,62,26,26,35,38,7,7,31,31,39,39,37,37,37,37,79,79,41,41,79,79,123,123,75,75,75),
(67,67,67,32,32,15,42,69,47,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,48,62,62,62,62,62,62,62,62,62,62,62,26,26,35,35,7,7,45,31,39,39,37,37,37,37,79,79,41,41,79,79,123,123,75,75,75),
(67,67,67,32,32,42,42,47,47,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,48,48,48,48,48,48,48,48,48,48,48,48,62,62,38,1,45,45,51,51,39,75,37,37,37,37,41,41,79,79,37,37,103,103,75,75,75),
(67,67,67,32,32,42,15,47,47,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,2,48,48,48,48,48,48,48,48,48,48,48,48,62,62,38,126,45,45,51,51,75,75,37,37,37,37,41,41,79,79,37,37,103,103,75,75,75),
(67,67,67,32,32,42,42,47,47,49,49,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,16,16,16,16,16,16,16,16,16,16,16,26,26,1,1,45,45,51,51,123,103,37,37,79,79,41,41,79,79,37,37,75,75,75,75,75),
(67,67,67,32,32,42,42,54,54,49,49,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,2,16,16,16,16,16,16,16,16,16,16,16,16,26,26,1,30,45,45,51,51,123,123,37,37,79,79,41,41,79,79,37,37,75,75,75,75,75),
(67,67,67,119,119,42,42,54,54,29,29,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,48,48,48,48,48,48,48,48,48,48,48,48,48,48,48,48,26,26,1,126,45,45,51,51,123,123,37,37,79,79,41,41,79,79,37,37,75,75,75,75,75),
(67,67,67,119,119,42,32,54,54,29,29,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,48,48,48,48,48,48,48,48,48,48,48,48,48,48,48,48,26,26,1,7,45,45,51,51,75,123,37,37,79,79,41,41,79,79,37,37,75,75,75,75,75),
(67,67,67,119,119,32,32,15,15,69,47,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,48,48,48,48,48,48,48,48,48,48,48,48,48,48,48,48,48,48,62,62,38,38,45,45,51,51,39,75,37,37,79,79,41,41,79,79,37,37,103,103,75,75,75),
(67,67,67,119,119,32,32,15,15,47,69,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,48,48,48,48,48,48,48,48,48,48,48,48,48,48,48,48,48,48,62,62,38,126,45,45,51,51,75,75,37,37,79,79,41,41,79,79,37,37,103,103,75,75,75),
(67,67,67,67,67,32,32,42,42,54,54,29,29,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,48,48,48,48,48,48,62,62,62,62,62,62,62,62,62,62,62,62,62,62,26,26,38,35,7,30,31,31,39,39,79,79,79,79,36,36,41,41,79,79,123,123,75,75,75),
(67,67,67,67,67,32,32,42,42,54,54,29,29,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,2,48,48,48,48,48,48,62,62,62,62,62,62,62,62,62,62,62,62,62,62,26,26,35,126,7,7,31,31,39,39,46,79,79,79,36,36,41,41,79,79,123,123,75,75,75),
(67,67,67,67,67,119,119,32,32,15,15,69,47,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,48,48,48,48,62,62,62,62,26,26,26,26,35,35,35,35,35,35,35,35,35,35,35,1,7,7,31,31,39,39,36,79,36,36,41,41,41,41,79,79,37,37,103,103,75),
(67,67,67,67,67,119,119,32,32,15,15,47,69,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,2,48,48,48,48,62,62,62,62,26,26,26,26,35,35,35,35,35,35,35,35,35,35,30,35,7,7,31,45,39,39,46,79,36,36,41,41,41,41,79,79,37,37,103,103,75),
(67,67,67,67,67,67,67,32,32,42,42,54,54,29,29,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,48,48,48,48,48,48,62,62,26,26,22,22,22,22,22,22,22,22,22,22,22,22,22,22,22,3,61,61,59,59,33,33,41,41,41,41,36,36,36,36,41,41,37,37,123,123,75),
(67,67,67,67,67,67,67,32,32,42,42,54,54,29,29,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,48,48,48,48,48,48,62,62,26,26,22,22,22,22,22,22,22,22,22,22,22,22,22,22,3,22,61,61,59,59,33,33,41,33,41,41,36,36,36,36,41,41,37,37,123,123,75),
(67,67,67,67,67,67,67,119,119,32,32,42,15,54,54,29,29,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,48,48,62,62,62,62,26,26,35,35,22,22,30,30,23,23,20,23,30,30,20,23,23,23,30,7,3,3,59,59,31,33,33,41,41,41,36,36,79,79,41,41,79,79,37,37,103),
(67,67,67,67,67,67,67,119,119,32,32,15,42,54,47,29,29,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,48,48,62,62,62,62,26,26,35,35,22,22,30,30,23,23,23,20,30,30,23,20,23,23,7,30,3,3,59,61,33,31,41,33,41,41,36,36,79,79,41,41,37,79,37,37,103),
(67,67,67,67,67,67,67,67,67,119,119,32,32,15,15,54,54,29,29,16,16,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,48,48,62,62,26,26,35,35,35,35,22,22,30,30,1,1,1,1,1,1,1,1,1,38,1,30,7,7,7,25,25,20,33,33,46,46,79,79,37,37,37,37,41,41,37,37,103),
(67,67,67,67,67,67,67,67,67,119,119,32,32,15,42,47,47,69,29,16,16,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,48,48,62,62,26,26,35,35,35,35,3,3,30,30,1,1,1,1,1,1,1,1,1,1,1,1,30,30,25,25,20,25,41,33,81,81,79,79,37,37,37,37,41,41,37,37,103),
(67,67,67,67,67,67,67,67,67,67,67,119,119,32,32,42,15,54,54,69,47,29,29,16,16,16,16,2,2,2,2,2,2,2,2,2,2,62,48,26,26,22,22,22,22,3,3,22,22,30,30,20,20,20,20,38,38,20,20,20,20,1,1,3,3,61,3,25,25,33,33,76,81,37,37,123,123,123,123,37,37,123,123,103),
(67,67,67,67,67,67,67,67,67,67,67,119,119,32,32,15,42,54,54,47,69,29,29,16,16,16,16,2,2,2,2,2,2,2,2,2,2,48,62,26,26,22,22,22,22,22,22,3,3,30,30,20,20,20,20,38,38,20,20,20,20,1,1,22,22,61,61,20,25,33,33,76,81,37,37,123,123,123,123,37,37,123,123,103),
(67,67,67,67,67,67,67,67,67,67,67,67,67,119,119,32,32,42,42,15,15,54,54,69,69,16,16,16,16,2,2,2,2,2,2,2,2,62,48,26,26,22,22,30,30,7,30,3,22,1,1,1,1,38,38,38,38,1,1,1,1,1,1,7,7,25,25,45,31,51,51,123,75,103,103,75,75,103,103,103,103,103,103,75),
(67,67,67,67,67,67,67,67,67,67,67,67,67,119,119,32,32,42,42,15,15,47,54,49,69,16,16,16,16,2,2,2,2,2,2,2,2,48,62,26,26,22,22,30,30,30,30,3,3,1,1,1,1,38,38,38,38,38,1,1,1,30,1,7,7,25,7,31,45,51,51,123,123,103,103,75,75,103,103,103,103,103,103,75),
(67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,119,119,32,32,32,32,42,42,15,15,16,29,16,16,2,2,2,2,2,2,2,2,16,16,29,29,22,22,30,30,23,23,22,22,30,30,20,20,20,20,30,30,23,23,23,23,30,7,3,61,59,59,33,33,39,39,103,123,75,75,75,75,75,75,75,75,75,75,75),
(67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,119,119,32,32,32,32,42,15,15,15,16,29,16,16,2,2,2,2,2,2,2,2,16,16,29,29,22,22,30,30,23,23,3,3,30,30,20,20,20,20,30,30,23,20,23,23,7,30,61,61,59,59,33,33,39,39,103,123,75,75,75,75,75,75,75,75,75,75,75),
(67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,119,119,32,32,15,15,29,69,16,16,2,2,2,2,2,2,2,2,16,16,29,29,22,22,30,30,30,30,22,22,30,30,30,30,30,30,22,3,22,3,3,3,3,3,61,61,59,59,33,33,79,46,37,37,75,75,75,75,75,75,75,75,75,75,75),
(67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,119,119,32,32,15,15,69,69,16,16,2,2,2,2,2,2,2,2,16,16,29,29,22,22,30,30,30,30,3,3,30,30,30,30,30,30,3,22,3,22,3,3,3,3,61,61,59,59,33,33,46,46,37,37,75,75,75,75,75,75,75,75,75,75,75),
(67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,119,119,32,32,15,15,69,69,16,16,2,2,2,2,2,2,2,2,16,16,29,29,22,22,30,30,7,7,3,3,60,60,60,60,60,60,3,3,7,7,30,30,7,7,25,25,31,33,33,41,46,46,37,37,103,103,75,75,75,75,75,75,75,75,75),
(67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,119,119,32,32,15,15,69,69,16,16,2,2,2,2,2,2,2,2,16,16,29,29,22,22,30,30,30,30,3,3,60,60,60,60,60,60,3,3,30,30,30,30,7,7,25,25,31,31,33,41,46,46,37,37,103,103,75,75,75,75,75,75,75,75,75),
(67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,32,32,42,42,54,54,29,29,16,16,2,2,2,2,2,2,2,2,16,16,29,29,22,22,23,60,60,60,3,3,60,60,60,60,60,60,3,3,7,7,23,23,24,24,25,25,31,31,81,46,41,41,37,37,123,123,75,75,75,75,75,75,75,75,75),
(67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,32,32,42,42,54,54,29,29,16,16,2,2,2,2,2,2,2,2,16,16,29,29,22,22,23,23,60,60,3,3,60,60,60,60,60,60,3,3,7,30,60,23,24,24,25,25,33,33,81,39,41,41,37,37,123,123,75,75,75,75,75,75,75,75,75),
(67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,119,119,32,32,15,15,69,69,16,16,2,2,2,2,2,2,2,2,2,2,16,16,29,29,22,22,3,3,3,3,3,3,3,3,3,3,3,3,3,3,30,7,7,7,25,7,45,45,51,51,46,79,41,41,79,79,37,37,103,103,103,103,103,103,103,103,75),
(67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,119,119,32,32,15,15,47,47,16,16,2,2,2,2,2,2,2,2,2,2,16,16,29,29,22,22,3,3,3,3,3,3,3,3,3,61,3,61,3,61,7,7,7,7,25,25,45,45,51,51,46,46,41,41,79,79,37,37,103,103,103,103,103,103,103,103,75),
(67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,119,119,42,42,54,54,29,29,16,16,2,2,2,2,2,2,16,16,16,16,29,29,29,29,69,47,47,47,47,47,47,47,54,54,30,30,60,60,3,3,60,60,60,60,18,18,31,31,39,39,79,79,79,79,41,41,79,79,37,37,37,37,37,37,123,123,103),
(67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,119,119,42,32,54,54,29,29,16,16,2,2,2,2,2,2,16,16,16,16,49,29,29,29,47,69,47,47,47,47,47,47,47,54,30,35,60,60,3,3,60,60,24,60,18,18,31,31,39,39,79,79,79,79,41,41,79,79,37,37,37,37,37,37,123,123,103),
(67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,32,32,42,42,47,47,49,49,2,2,2,2,2,2,16,16,16,16,29,29,22,22,22,22,22,22,22,22,22,22,22,22,3,22,3,3,3,3,3,3,3,3,3,61,61,59,31,33,39,39,46,79,37,37,41,41,79,79,79,79,79,79,41,41,37,37,103),
(67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,32,32,42,42,47,54,49,49,2,2,2,2,2,2,16,16,16,16,49,29,22,22,22,22,22,22,22,22,22,22,22,22,22,3,3,3,3,3,3,3,3,3,61,61,59,59,31,31,39,39,79,79,37,37,41,41,79,79,79,79,79,79,41,41,37,37,103),
(67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,32,32,42,42,69,47,16,16,2,2,2,2,2,2,16,16,20,20,20,20,22,22,30,30,30,30,1,1,1,1,1,1,1,38,1,1,1,30,30,30,30,30,7,7,7,25,31,31,39,39,81,81,37,37,79,79,41,41,41,41,41,41,79,79,37,37,103),
(67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,32,32,15,42,69,47,16,16,2,2,2,2,2,2,16,16,20,20,20,20,22,22,30,30,1,30,1,1,1,1,1,1,1,1,1,1,1,1,30,30,30,30,7,7,25,25,45,45,39,51,81,81,37,37,79,79,41,41,41,41,41,41,79,79,37,37,103),
(67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,32,32,42,42,47,47,16,16,2,2,2,2,16,16,16,16,20,20,30,30,3,3,30,30,23,20,20,20,1,1,20,20,20,20,38,38,38,38,20,20,20,20,1,1,24,60,59,59,31,33,39,39,123,123,37,37,79,79,36,36,41,41,79,79,123,123,75),
(67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,32,32,42,15,47,47,16,16,2,2,2,2,16,16,16,16,20,20,30,30,3,3,30,30,20,23,20,20,1,1,20,20,20,20,38,38,38,38,20,20,20,20,1,1,24,24,59,59,33,31,39,81,123,123,37,37,79,79,36,36,41,41,79,79,123,123,75),
(67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,32,32,42,42,47,47,49,49,2,2,2,2,16,16,49,49,20,20,30,30,22,3,1,1,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,7,7,25,25,45,45,39,51,123,123,37,37,79,79,41,41,79,79,37,37,103,103,75),
(67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,32,32,42,42,54,54,49,49,2,2,2,2,16,16,49,49,20,20,30,30,3,22,1,1,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,1,1,25,25,31,45,51,51,123,123,37,37,79,79,41,41,79,79,37,37,103,103,75),
(67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,119,119,42,42,54,54,29,29,16,16,2,2,16,16,29,29,22,22,22,22,22,3,1,1,20,20,20,20,38,38,20,20,20,20,38,38,38,38,20,20,20,20,38,38,23,20,3,3,25,25,41,33,81,81,79,79,79,79,41,41,37,37,123,123,75,75,75),
(67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,119,119,42,32,54,54,29,29,16,16,2,2,16,16,29,29,22,22,22,22,3,22,1,1,20,20,20,20,38,38,20,20,20,20,38,38,38,38,20,25,20,20,38,38,20,23,61,61,25,25,33,33,76,81,79,79,36,79,41,41,37,37,123,123,75,75,75),
(67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,119,119,32,32,15,15,47,47,16,16,2,2,16,16,29,29,22,22,30,30,1,30,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,1,38,7,7,25,25,41,33,76,81,36,36,41,41,79,79,37,37,103,103,75,75,75),
(67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,119,119,32,32,15,15,69,69,16,16,2,2,16,16,29,29,22,22,30,30,30,1,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,1,1,7,7,25,25,33,33,76,81,36,36,41,41,79,79,37,37,103,103,75,75,75),
(67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,32,32,42,42,54,54,29,29,16,16,16,16,29,29,22,22,30,30,20,23,1,1,20,20,20,20,1,1,20,20,20,20,38,38,38,38,20,20,20,20,1,1,23,23,61,61,45,31,51,39,41,41,41,41,41,41,79,79,37,37,75,75,75,75,75),
(67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,32,32,42,42,54,54,29,29,16,16,16,16,29,29,22,22,30,30,23,20,1,1,20,20,20,20,1,1,20,20,20,20,38,38,38,38,20,20,20,20,1,1,23,24,61,61,31,45,39,51,41,41,41,41,41,41,79,79,37,37,75,75,75,75,75),
(67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,119,119,32,32,15,15,69,69,16,16,16,16,49,49,22,22,1,30,30,30,1,1,30,30,30,30,30,30,30,30,30,30,1,1,1,1,30,30,30,30,30,30,7,7,25,25,31,33,39,39,36,36,36,36,41,41,79,79,37,37,75,75,75,75,75),
(67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,119,119,32,32,15,15,69,69,16,16,16,16,49,49,22,22,38,1,30,30,1,1,30,30,30,30,30,30,30,30,30,30,30,1,30,1,30,30,30,30,7,7,7,7,25,25,33,31,39,81,36,36,36,36,41,41,79,79,37,37,75,75,75,75,75),
(67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,119,119,32,32,15,15,69,69,16,16,16,16,49,49,22,22,22,22,22,22,22,22,3,3,3,3,3,3,3,3,3,3,22,3,22,3,22,3,3,3,3,3,61,59,45,31,51,39,46,46,36,36,41,41,41,41,36,36,37,37,103,103,75,75,75),
(67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,119,119,32,32,15,15,29,69,16,16,16,16,49,49,22,22,22,22,22,22,22,22,3,3,3,3,3,3,3,3,3,3,3,22,3,22,3,22,3,3,3,3,61,61,31,45,39,51,46,79,36,36,41,41,41,41,36,36,37,37,103,103,75,75,75),
(67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,119,119,32,32,42,42,15,15,69,29,16,16,2,2,16,16,49,2,49,16,29,29,69,69,3,3,60,60,3,3,60,60,23,23,23,23,23,23,23,23,23,23,60,24,18,18,31,31,39,39,79,79,79,79,41,41,36,36,41,41,37,37,123,123,75,75,75),
(67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,119,119,32,32,42,42,15,59,69,29,16,16,2,2,16,16,49,49,49,49,29,29,69,69,3,3,60,60,3,3,60,60,23,23,23,23,23,23,23,23,23,23,24,60,18,18,31,31,39,39,79,79,79,79,41,41,36,36,41,41,37,37,123,123,75,75,75),
(67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,119,119,32,32,42,15,54,54,69,47,16,16,16,16,2,2,2,2,16,16,16,16,49,49,29,29,22,22,30,7,3,3,30,30,30,30,1,1,1,1,1,1,1,1,7,7,25,25,31,31,39,39,79,79,41,41,36,36,36,36,41,41,79,79,37,37,123,123,75),
(67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,119,119,32,32,15,42,54,54,69,69,16,16,16,16,2,2,2,2,16,16,16,16,49,49,29,29,22,3,30,7,3,3,30,30,30,30,38,1,1,1,1,1,1,1,7,7,25,25,31,31,39,39,79,79,41,41,36,36,36,36,41,41,79,79,37,37,123,123,75),
(67,67,67,67,67,67,67,67,67,67,67,67,67,119,119,32,32,15,15,54,47,29,29,16,16,16,16,2,2,2,2,2,2,2,2,2,2,16,16,49,49,22,22,22,3,3,22,30,30,1,1,20,20,20,20,38,38,20,20,20,20,7,7,45,45,51,51,79,46,41,41,79,79,36,36,36,36,41,41,79,79,37,37,103),
(67,67,67,67,67,67,67,67,67,67,67,67,67,119,119,32,32,15,42,47,54,29,29,16,16,16,16,2,2,2,2,2,2,2,2,2,2,16,16,49,49,22,22,22,22,22,3,30,1,1,1,20,20,20,20,38,38,20,20,20,20,25,7,45,45,51,51,46,46,41,41,79,79,36,36,36,36,41,41,79,79,37,37,103),
(67,67,67,67,67,67,67,67,67,67,67,119,119,32,32,42,15,54,47,29,29,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,29,49,69,69,22,22,1,1,38,38,38,38,38,38,38,38,38,38,38,38,7,7,25,25,31,31,76,81,41,41,36,36,36,36,36,36,41,41,41,41,37,37,103),
(67,67,67,67,67,67,67,67,67,67,67,119,119,32,32,15,42,47,54,29,29,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,29,29,69,69,22,22,1,1,38,38,38,38,38,38,38,38,38,38,38,38,7,7,25,25,31,31,39,76,41,41,36,36,36,36,36,36,41,41,41,41,37,37,103),
(67,67,67,67,67,67,67,67,67,67,67,32,32,42,42,54,54,29,29,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,29,29,22,22,1,1,1,1,20,20,20,20,1,1,20,20,20,20,1,7,24,24,45,31,39,39,41,41,36,36,41,41,41,41,79,79,37,37,123,123,103),
(67,67,67,67,67,67,67,67,67,67,67,32,32,42,42,54,54,29,29,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,29,29,22,22,1,1,1,1,20,20,20,20,1,1,20,20,20,20,7,1,18,24,31,45,39,39,41,41,36,36,41,41,41,41,79,79,37,37,123,123,103),
(67,67,67,67,67,67,67,67,67,119,119,32,32,15,15,69,47,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,29,29,22,22,30,30,30,30,1,1,1,1,1,1,1,1,1,1,30,30,7,7,25,25,33,33,46,46,41,41,79,79,79,79,37,37,123,123,103,103,75),
(67,67,67,67,67,67,67,67,67,119,119,32,32,15,15,47,69,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,29,29,22,22,38,1,30,30,38,1,1,1,1,1,1,1,1,1,30,30,7,7,25,25,33,33,81,46,41,41,79,79,79,79,37,37,123,123,103,103,75),
(67,67,67,67,67,67,67,67,67,32,32,42,42,54,54,29,29,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,49,49,22,22,22,22,22,22,22,22,22,22,22,22,22,22,22,22,22,22,22,3,61,61,31,31,39,39,41,41,79,79,37,37,103,103,75,75,75,75,75),
(67,67,67,67,67,67,67,67,67,32,32,42,42,54,54,29,29,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,49,49,22,22,22,22,22,22,22,22,22,22,22,22,22,22,22,22,22,22,3,3,61,61,31,31,39,39,41,41,79,79,37,37,103,103,75,75,75,75,75),
(67,67,67,67,67,67,67,119,119,32,32,15,15,69,47,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,49,16,62,62,26,26,26,26,26,26,26,26,26,26,26,26,26,26,35,35,30,30,59,59,33,33,81,81,37,37,103,103,75,75,75,75,75,75,75),
(67,67,67,67,67,67,67,119,119,32,32,15,15,47,69,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,49,16,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,35,35,30,126,59,59,33,33,81,81,37,37,103,103,75,75,75,75,75,75,75),
(67,67,67,67,67,67,67,119,119,42,42,54,54,29,29,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,62,48,62,62,62,62,62,62,62,62,62,62,62,62,62,62,26,26,1,38,25,25,33,33,76,81,123,123,75,75,75,75,75,75,75,75,75),
(67,67,67,67,67,67,67,119,119,42,32,54,54,29,29,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,48,62,62,62,62,62,62,62,62,62,62,62,62,62,62,62,26,26,126,30,7,7,31,31,81,81,123,123,75,75,75,75,75,75,75,75,75),
(67,67,67,67,67,67,67,32,32,42,42,47,47,49,49,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,16,16,16,16,16,16,16,16,16,16,16,48,48,48,48,26,26,38,38,45,45,51,51,75,75,103,103,75,75,75,75,75,75,75,75,75),
(67,67,67,67,67,67,67,32,32,42,42,47,54,49,49,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,2,16,16,16,16,16,16,16,16,16,16,16,16,48,48,48,48,26,26,38,126,45,45,51,51,75,75,103,103,75,75,75,75,75,75,75,75,75),
(67,67,67,67,67,67,67,32,32,42,42,69,47,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,48,48,48,48,48,48,48,48,48,48,48,48,48,48,48,48,48,48,48,48,26,26,7,1,45,45,39,51,123,103,75,75,75,75,75,75,75,75,75,75,75),
(67,67,67,67,67,67,67,32,32,15,42,69,47,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,48,48,48,48,48,48,48,48,48,48,48,48,48,48,48,48,48,48,62,48,26,26,1,7,45,45,51,39,123,123,75,75,75,75,75,75,75,75,75,75,75),
(67,67,67,67,67,67,67,32,32,42,42,47,47,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,48,48,48,48,48,48,48,48,48,48,48,48,48,48,48,48,48,48,48,48,62,62,38,38,7,7,31,33,76,39,37,37,75,75,75,75,75,75,75,75,75,75,75),
(67,67,67,67,67,67,67,32,32,42,15,47,47,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,48,48,48,48,48,48,48,48,48,48,48,48,48,48,48,48,48,48,48,48,62,62,35,26,7,7,31,31,76,76,37,37,75,75,75,75,75,75,75,75,75,75,75),
(67,67,67,67,67,67,67,32,32,42,42,47,47,49,49,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,48,48,48,48,48,48,62,62,62,62,62,62,62,62,62,62,62,62,62,62,62,62,26,26,1,7,45,45,33,33,76,76,37,37,103,103,75,75,75,75,75,75,75,75,75),
(67,67,67,67,67,67,67,32,32,42,42,54,54,49,49,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,2,48,48,48,48,48,48,62,62,62,62,62,62,62,62,62,62,62,62,62,62,62,62,26,26,30,1,45,45,33,33,76,76,37,37,103,103,75,75,75,75,75,75,75,75,75),
(67,67,67,67,67,67,67,119,119,42,42,54,54,29,29,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,48,48,48,48,62,62,62,62,26,26,26,26,35,35,35,35,35,35,35,35,35,35,30,38,7,7,31,31,39,76,41,41,37,37,123,123,75,75,75,75,75,75,75,75,75),
(67,67,67,67,67,67,67,119,119,42,32,54,54,29,29,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,2,48,48,48,48,62,62,62,62,26,26,26,26,35,35,35,35,35,35,35,35,35,35,35,35,7,7,31,31,39,39,41,41,37,37,123,123,75,75,75,75,75,75,75,75,75),
(67,67,67,67,67,67,67,119,119,32,32,15,15,69,47,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,48,48,48,48,48,48,62,62,26,26,22,22,22,22,22,22,22,22,22,22,22,22,22,3,61,61,45,45,51,51,46,79,41,41,79,79,37,37,103,103,75,75,75,75,75,75,75),
(67,67,67,67,67,67,67,119,119,32,32,15,15,47,69,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,48,48,48,48,48,48,62,62,26,26,22,22,22,22,22,22,22,22,22,22,22,22,3,3,61,61,45,45,51,51,46,46,41,41,79,79,37,37,103,103,75,75,75,75,75,75,75),
(67,67,67,67,67,67,67,67,67,32,32,42,42,54,54,29,29,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,48,48,62,62,62,62,26,26,35,35,22,22,30,30,23,23,20,23,30,30,20,23,23,23,25,25,45,31,51,39,79,79,79,79,41,41,79,79,37,37,103,103,75,75,75,75,75),
(67,67,67,67,67,67,67,67,67,32,32,42,42,54,54,29,29,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,48,48,62,62,62,62,26,26,35,35,22,22,30,30,23,23,23,20,30,30,23,20,23,24,25,25,31,31,39,51,79,79,79,79,41,41,79,79,37,37,103,103,75,75,75,75,75),
(67,67,67,67,67,67,67,67,67,119,119,32,32,15,15,69,47,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,48,48,62,62,26,26,35,35,35,35,22,22,30,30,1,1,1,1,1,1,1,1,7,7,25,7,45,45,39,39,79,79,37,37,41,41,79,79,79,79,37,37,123,123,103,103,75),
(67,67,67,67,67,67,67,67,67,119,119,32,32,15,15,47,69,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,48,48,62,62,26,26,35,35,35,35,3,3,30,30,1,1,1,1,1,1,1,1,7,7,25,25,45,31,51,39,79,79,37,37,41,41,79,79,79,79,37,37,123,123,103,103,75),
(67,67,67,67,67,67,67,67,67,67,67,32,32,42,42,54,54,29,29,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,62,48,26,26,22,22,22,22,3,3,22,22,30,30,20,20,20,20,38,38,20,20,20,20,7,7,45,45,51,51,76,76,37,37,79,79,41,41,41,41,79,79,37,37,123,123,103),
(67,67,67,67,67,67,67,67,67,67,67,32,32,42,42,54,54,69,29,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,48,62,26,26,22,22,22,22,22,22,3,3,30,30,20,20,20,20,38,38,20,20,20,20,25,7,45,45,51,51,76,76,37,37,79,79,41,41,41,41,79,79,37,37,123,123,103),
(67,67,67,67,67,67,67,67,67,67,67,119,119,32,32,42,15,47,54,29,29,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,62,48,26,26,22,22,30,30,7,30,3,22,1,1,1,1,38,38,38,38,1,1,1,1,7,7,25,25,33,31,76,81,37,37,37,37,79,79,36,36,41,41,41,41,37,37,103),
(67,67,67,67,67,67,67,67,67,67,67,119,119,32,32,15,42,54,47,29,29,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,48,62,26,26,22,22,30,30,30,30,3,3,1,1,1,1,38,38,38,38,38,1,1,1,7,7,25,25,33,33,81,81,37,37,37,37,79,79,36,36,41,41,41,41,37,37,103),
(67,67,67,67,67,67,67,67,67,67,67,67,67,119,119,32,32,15,15,54,47,49,49,16,16,2,2,2,2,2,2,2,2,2,2,2,2,16,16,29,29,22,22,30,30,23,23,22,22,30,30,20,20,20,20,30,30,23,23,23,23,7,7,18,18,33,31,81,81,37,37,37,37,37,37,36,36,41,41,79,79,37,37,103),
(67,67,67,67,67,67,67,67,67,67,67,67,67,119,119,32,32,15,15,69,47,16,49,16,16,2,2,2,2,2,2,2,2,2,2,2,2,16,16,29,29,22,22,30,30,23,23,3,3,30,30,20,20,20,20,30,30,23,20,23,23,7,7,18,18,33,33,81,81,37,37,37,37,37,37,36,36,41,41,79,79,37,37,103),
(67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,119,119,42,32,15,15,16,29,16,16,2,2,2,2,2,2,2,2,2,2,2,2,16,16,29,29,22,22,30,30,30,30,22,22,30,30,30,30,30,30,22,3,22,3,3,3,61,61,59,59,33,33,41,41,79,79,79,79,79,79,41,41,79,79,37,37,123,123,75),
(67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,119,119,32,42,15,15,16,29,16,16,2,2,2,2,2,2,2,2,2,2,2,2,16,16,29,29,22,22,30,30,30,30,3,3,30,30,30,30,30,30,3,22,3,22,3,3,61,3,59,59,33,33,41,41,79,79,79,79,79,79,41,41,79,79,37,37,123,123,75),
(67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,119,119,42,42,15,15,16,29,16,16,2,2,2,2,2,2,2,2,2,2,2,2,16,16,29,29,22,22,30,30,7,7,3,3,60,60,60,60,60,60,3,3,7,7,7,30,7,7,20,25,33,33,41,41,79,79,36,36,36,36,41,41,37,37,123,123,75,75,75),
(67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,119,119,32,42,15,15,29,29,16,16,2,2,2,2,2,2,2,2,2,2,2,2,16,16,29,29,22,22,30,30,30,30,3,3,60,60,60,60,60,60,3,3,30,30,7,7,7,25,25,25,33,33,41,41,36,36,36,36,36,36,41,41,37,37,123,123,75,75,75),
(67,67,67,67,67,67,67,67,67,67,67,67,67,119,119,32,32,15,15,47,47,49,49,16,16,2,2,2,2,2,2,2,2,2,2,2,2,16,16,29,29,22,22,23,60,60,60,3,3,60,60,60,60,60,60,3,3,7,7,23,23,18,24,31,31,51,39,46,46,41,41,41,41,41,41,79,79,37,37,103,103,75,75,75),
(67,67,67,67,67,67,67,67,67,67,67,67,67,119,119,32,32,15,42,47,47,49,49,16,16,2,2,2,2,2,2,2,2,2,2,2,2,16,16,29,29,22,22,23,23,60,60,3,3,60,60,60,60,60,60,3,3,7,30,60,23,24,24,45,45,39,39,46,46,41,41,41,41,41,41,79,79,37,37,103,103,75,75,75),
(67,67,67,67,67,67,67,67,67,67,67,67,67,32,32,42,42,54,54,29,29,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,29,29,22,22,3,3,3,3,3,3,3,3,3,3,3,3,3,3,30,7,7,7,25,25,31,31,39,39,79,79,79,79,36,36,41,41,79,79,37,37,75,75,75,75,75),
(67,67,67,67,67,67,67,67,67,67,67,67,67,32,32,42,42,54,54,29,29,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,29,29,22,22,3,3,3,3,3,3,3,3,3,61,3,61,3,61,7,7,7,7,25,25,31,31,39,39,79,79,79,79,36,36,41,41,79,79,37,37,75,75,75,75,75),
(67,67,67,67,67,67,67,67,67,67,67,119,119,32,32,15,15,69,47,16,16,2,2,2,2,2,2,2,2,2,2,2,2,16,16,16,16,29,29,29,29,69,47,47,47,47,47,47,47,54,54,30,30,60,60,3,3,60,60,60,18,18,18,31,31,39,39,37,37,79,79,36,36,41,41,79,79,37,37,75,75,75,75,75),
(67,67,67,67,67,67,67,67,67,67,67,119,119,32,32,15,15,47,69,16,16,2,2,2,2,2,2,2,2,2,2,2,2,16,16,16,16,49,29,29,29,47,69,47,47,47,47,47,47,47,54,30,35,60,60,3,3,60,60,24,60,18,18,31,31,39,39,37,37,79,79,36,36,41,41,79,79,37,37,75,75,75,75,75),
(67,67,67,67,67,67,67,67,67,67,67,32,32,42,42,54,54,29,29,16,16,2,2,2,2,2,2,2,2,2,2,16,16,16,16,29,29,22,22,22,22,22,22,22,22,22,22,22,22,3,22,3,3,3,3,3,3,3,3,3,3,61,61,45,45,39,51,76,76,79,79,41,41,41,41,36,36,37,37,103,103,75,75,75),
(67,67,67,67,67,67,67,67,67,67,67,32,32,42,42,54,54,29,29,16,16,2,2,2,2,2,2,2,2,2,2,16,16,16,16,49,29,22,22,22,22,22,22,22,22,22,22,22,22,22,3,3,3,3,3,3,3,3,3,3,3,61,61,45,31,51,51,76,76,79,79,41,41,41,41,36,36,37,37,103,103,75,75,75),
(67,67,67,67,67,67,67,67,67,119,119,32,32,15,15,69,47,16,16,2,2,2,2,2,2,2,2,2,2,2,2,16,16,20,20,20,20,22,22,30,30,30,30,1,1,1,1,1,1,1,38,1,1,1,30,30,30,30,30,7,7,7,7,25,25,33,31,39,39,36,36,41,41,36,36,41,41,37,37,123,123,75,75,75),
(67,67,67,67,67,67,67,67,67,119,119,32,32,15,15,47,69,16,16,2,2,2,2,2,2,2,2,2,2,2,2,16,16,20,20,20,20,22,22,30,30,1,30,1,1,1,1,1,1,1,1,1,1,1,1,30,30,30,30,30,30,7,7,25,25,31,31,76,39,36,36,41,41,36,36,41,41,37,37,123,123,75,75,75),
(67,67,67,67,67,67,67,67,67,119,119,42,42,54,54,29,29,16,16,2,2,2,2,2,2,2,2,2,2,16,16,16,16,20,20,30,30,3,3,30,30,23,20,20,20,1,1,20,20,20,20,38,38,38,38,20,20,20,20,1,1,23,24,24,18,45,31,51,39,41,41,36,36,36,36,41,41,79,79,37,37,103,103,75),
(67,67,67,67,67,67,67,67,67,119,119,42,32,54,54,29,29,16,16,2,2,2,2,2,2,2,2,2,2,16,16,16,16,20,20,30,30,3,3,30,30,20,23,20,20,1,1,20,20,20,20,38,38,38,38,20,20,20,20,1,1,23,20,24,24,45,45,51,51,41,41,36,36,36,36,41,41,79,79,37,37,103,103,75),
(67,67,67,67,67,67,67,67,67,32,32,42,42,47,47,49,49,2,2,2,2,2,2,2,2,2,2,2,2,16,16,49,49,20,20,30,30,22,3,1,1,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,1,7,7,25,25,33,33,41,41,79,36,79,79,79,79,41,41,37,37,123,123,75),
(67,67,67,67,67,67,67,67,67,32,32,42,42,47,54,49,49,2,2,2,2,2,2,2,2,2,2,2,2,16,16,49,49,20,20,30,30,3,22,1,1,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,7,7,25,25,31,31,41,41,36,36,79,79,79,79,41,41,37,37,123,123,75),
(67,67,67,67,67,67,67,67,67,32,32,42,42,69,47,16,16,2,2,2,2,2,2,2,2,2,2,2,2,16,16,29,29,22,22,22,22,22,3,1,1,20,20,20,20,38,38,20,20,20,20,38,38,38,38,20,20,20,20,38,38,20,20,20,20,25,25,45,45,33,33,46,79,37,37,37,37,41,41,79,79,37,37,103),
(67,67,67,67,67,67,67,67,67,32,32,15,42,69,47,16,16,2,2,2,2,2,2,2,2,2,2,2,2,16,16,29,29,22,22,22,22,3,22,1,1,20,20,20,20,38,38,20,20,20,20,38,38,38,38,20,25,20,20,38,38,20,20,20,20,25,7,31,31,41,41,46,79,37,37,37,37,41,41,37,79,37,37,103),
(67,67,67,67,67,67,67,67,67,32,32,42,42,47,47,16,16,2,2,2,2,2,2,2,2,2,2,2,2,16,16,29,29,22,22,30,30,1,30,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,1,1,7,7,25,25,33,33,76,81,37,37,37,37,37,37,41,41,37,37,103),
(67,67,67,67,67,67,67,67,67,32,32,42,15,47,47,16,16,2,2,2,2,2,2,2,2,2,2,2,2,16,16,29,29,22,22,30,30,30,1,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,1,1,7,7,25,25,33,33,76,81,37,37,37,37,37,37,41,41,37,37,103),
(67,67,67,67,67,67,67,67,67,32,32,42,42,47,47,49,49,2,2,2,2,2,2,2,2,2,2,2,2,16,16,29,29,22,22,30,30,20,23,1,1,20,20,20,20,1,1,20,20,20,20,38,38,38,38,20,20,20,20,1,1,20,20,20,23,7,25,59,59,33,33,76,81,123,123,103,103,123,123,37,37,123,123,103),
(67,67,67,67,67,67,67,67,67,32,32,42,42,54,54,49,49,2,2,2,2,2,2,2,2,2,2,2,2,16,16,29,29,22,22,30,30,23,20,1,1,20,20,20,20,1,1,20,20,20,20,38,38,38,38,20,20,20,20,1,1,20,20,23,20,7,7,59,59,33,33,81,81,123,123,103,103,123,123,37,37,123,123,103),
(67,67,67,67,67,67,67,67,67,119,119,42,42,54,54,29,29,16,16,2,2,2,2,2,2,2,2,2,2,16,16,49,49,22,22,1,30,30,30,1,1,30,30,30,30,30,30,30,30,30,30,1,1,1,1,30,30,30,30,30,30,30,30,7,7,25,25,45,45,51,51,81,81,103,103,75,75,103,103,103,103,103,103,75),
(67,67,67,67,67,67,67,67,67,119,119,42,42,54,54,29,29,16,16,2,2,2,2,2,2,2,2,2,2,16,16,49,49,22,22,38,1,30,30,1,1,30,30,30,30,30,30,30,30,30,30,30,1,30,1,30,30,30,30,30,30,30,30,7,7,25,7,45,45,51,51,81,81,103,103,75,75,103,103,103,103,103,103,75),
(67,67,67,67,67,67,67,67,67,119,119,32,32,15,15,29,69,16,16,2,2,2,2,2,2,2,2,2,2,16,16,49,49,22,22,22,22,22,22,22,22,3,3,3,3,3,3,3,3,3,3,22,3,22,3,22,3,3,3,3,3,3,3,3,3,61,61,45,31,51,51,81,81,103,103,75,75,75,75,75,75,75,75,75),
(67,67,67,67,67,67,67,67,67,119,119,32,32,15,15,16,69,16,16,2,2,2,2,2,2,2,2,2,2,16,16,49,49,22,22,22,22,22,22,22,22,3,3,3,3,3,3,3,3,3,3,3,22,3,22,3,22,3,3,3,3,3,3,3,3,61,61,31,45,39,51,75,75,103,103,75,75,75,75,75,75,75,75,75),
(67,67,67,67,67,67,67,67,67,119,119,42,42,15,15,16,29,16,16,2,2,2,2,2,2,2,2,2,2,2,2,16,16,49,2,49,16,29,29,69,69,3,3,60,60,3,3,60,60,23,23,23,23,23,23,23,23,23,23,23,23,23,23,23,23,24,24,18,18,33,33,81,81,123,123,75,75,75,75,75,75,75,75,75),
(67,67,67,67,67,67,67,67,67,119,119,32,42,15,15,29,29,16,16,2,2,2,2,2,2,2,2,2,2,2,2,16,16,49,49,49,49,29,29,69,69,3,3,60,60,3,3,60,60,23,23,23,23,23,23,23,23,23,23,23,23,23,23,23,23,24,24,18,18,33,33,76,81,123,123,75,75,75,75,75,75,75,75,75),
(67,67,67,67,67,67,67,119,119,32,32,15,15,47,47,49,49,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,16,16,49,49,29,29,22,22,30,7,3,3,30,30,30,30,1,1,1,1,1,1,1,1,1,1,1,1,1,1,7,7,25,25,31,31,39,51,123,123,75,75,75,75,75,75,75,75,75),
(67,67,67,67,67,67,67,119,119,32,32,15,42,47,47,49,49,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,16,16,49,49,29,29,22,3,30,7,3,3,30,30,30,30,38,1,1,1,1,1,1,1,1,1,1,1,1,1,7,7,25,25,31,31,39,39,123,123,75,75,75,75,75,75,75,75,75),
(67,67,67,67,67,67,67,32,32,42,42,54,54,29,29,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,49,49,22,22,22,3,3,22,30,30,1,1,20,20,20,20,38,38,20,20,20,20,38,38,20,20,20,20,25,7,45,45,51,51,123,123,103,103,103,103,103,103,103,103,75),
(67,67,67,67,67,67,67,32,32,42,42,54,54,29,29,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,49,49,22,22,22,22,22,3,30,1,1,1,20,20,20,20,38,38,20,20,20,20,38,38,20,20,20,20,25,7,31,45,51,51,123,123,103,103,103,103,103,103,103,103,75),
(67,67,67,67,67,119,119,32,32,15,15,69,47,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,29,49,69,69,22,22,1,1,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,1,1,7,25,25,25,41,33,76,76,37,37,37,37,37,37,123,123,103),
(67,67,67,67,67,119,119,32,32,15,15,47,69,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,29,29,69,69,22,22,1,1,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,1,1,25,7,25,25,41,33,76,76,37,37,37,37,37,37,123,123,103),
(67,67,67,67,67,32,32,42,42,54,54,29,29,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,29,29,22,22,1,1,1,1,20,20,20,20,1,1,20,20,20,20,1,1,20,20,23,24,25,25,31,33,41,41,46,46,79,79,79,79,41,41,37,37,103),
(67,67,67,67,67,32,32,42,42,54,54,29,29,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,29,29,22,22,1,1,1,1,20,20,20,20,1,1,20,20,20,20,1,1,20,20,24,24,25,25,31,31,41,33,79,46,79,79,79,79,41,41,37,37,103),
(67,67,67,119,119,32,32,15,15,69,47,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,29,29,22,22,30,30,30,30,1,1,1,1,1,1,1,1,1,1,1,1,7,7,25,7,45,45,51,51,81,46,41,41,36,36,41,41,79,37,37,37,103),
(67,67,67,119,119,32,32,15,15,47,69,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,29,29,22,22,38,1,30,30,38,1,1,1,1,1,1,1,1,1,1,1,7,7,7,25,45,45,51,51,81,81,41,41,36,36,41,41,79,79,37,37,103),
(67,67,67,119,119,42,42,54,54,29,29,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,49,49,22,22,22,22,22,22,22,22,22,22,22,22,22,22,22,22,22,22,3,61,59,59,33,33,81,39,79,79,41,41,36,36,41,41,37,37,123,123,75),
(67,67,67,119,119,42,32,54,54,29,29,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,49,49,22,22,22,22,22,22,22,22,22,22,22,22,22,22,22,22,3,22,61,3,59,59,31,31,81,81,79,79,41,41,36,36,41,41,37,37,123,123,75),
(67,67,67,32,32,42,42,47,47,49,49,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,49,16,26,62,26,26,26,26,26,26,26,26,26,26,26,26,35,35,7,30,45,45,39,39,81,81,37,37,79,79,41,41,79,79,37,37,103,103,75),
(67,67,67,32,32,42,42,47,54,49,49,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,49,49,26,26,26,26,26,26,26,26,26,26,26,26,26,26,35,35,7,7,31,45,39,39,81,81,37,37,79,79,41,41,79,79,37,37,103,103,75),
(67,67,67,32,32,42,42,69,47,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,62,48,62,62,62,62,62,62,62,62,62,62,26,26,35,38,7,7,31,31,39,39,37,37,37,37,79,79,41,41,79,79,123,123,75,75,75),
(67,67,67,32,32,15,42,69,47,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,48,62,62,62,62,62,62,62,62,62,62,62,26,26,35,35,7,7,45,31,39,39,37,37,37,37,79,79,41,41,79,79,123,123,75,75,75),
(67,67,67,32,32,42,42,47,47,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,48,48,48,48,48,48,48,48,48,48,48,48,62,62,38,1,45,45,51,51,39,75,37,37,37,37,41,41,79,79,37,37,103,103,75,75,75),
(67,67,67,32,32,42,15,47,47,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,2,48,48,48,48,48,48,48,48,48,48,48,48,62,62,38,126,45,45,51,51,75,75,37,37,37,37,41,41,79,79,37,37,103,103,75,75,75),
(67,67,67,32,32,42,42,47,47,49,49,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,16,16,16,16,16,16,16,16,16,16,16,26,26,1,1,45,45,51,51,123,103,37,37,79,79,41,41,79,79,37,37,75,75,75,75,75),
(67,67,67,32,32,42,42,54,54,49,49,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,2,16,16,16,16,16,16,16,16,16,16,16,16,26,26,1,30,45,45,51,51,123,123,37,37,79,79,41,41,79,79,37,37,75,75,75,75,75),
(67,67,67,119,119,42,42,54,54,29,29,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,48,48,48,48,48,48,48,48,48,48,48,48,48,48,48,48,26,26,1,126,45,45,51,51,123,123,37,37,79,79,41,41,79,79,37,37,75,75,75,75,75),
(67,67,67,119,119,42,32,54,54,29,29,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,48,48,48,48,48,48,48,48,48,48,48,48,48,48,48,48,26,26,1,7,45,45,51,51,75,123,37,37,79,79,41,41,79,79,37,37,75,75,75,75,75),
(67,67,67,119,119,32,32,15,15,69,69,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,48,48,48,48,48,48,48,48,48,48,48,48,48,48,48,48,48,48,62,62,38,38,45,45,51,51,39,75,37,37,79,79,41,41,79,79,37,37,103,103,75,75,75),
(67,67,67,119,119,32,32,15,15,69,69,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,48,48,48,48,48,48,48,48,48,48,48,48,48,48,48,48,48,48,62,62,38,126,45,45,51,51,75,75,37,37,79,79,41,41,79,79,37,37,103,103,75,75,75),
(67,67,67,67,67,32,32,15,42,47,47,49,49,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,48,48,48,48,48,48,62,62,62,62,62,62,62,62,62,62,62,62,62,62,26,26,38,35,7,30,31,31,39,39,37,37,79,79,36,36,41,41,79,79,123,123,75,75,75),
(67,67,67,67,67,32,32,42,15,47,47,49,49,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,2,48,48,48,48,48,48,62,62,62,62,62,62,62,62,62,62,62,62,62,62,26,26,35,126,7,7,31,31,39,39,37,37,79,79,36,36,41,41,79,79,123,123,75,75,75),
(67,67,67,67,67,119,119,42,32,54,54,29,29,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,48,48,48,48,62,62,62,62,26,26,26,26,35,35,35,35,35,35,35,35,35,35,35,1,7,7,31,31,39,39,46,79,79,79,41,41,41,41,79,79,37,37,103,103,75),
(67,67,67,67,67,119,119,42,42,54,54,29,29,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,2,48,48,48,48,62,62,62,62,26,26,26,26,35,35,35,35,35,35,35,35,35,35,35,35,7,7,45,45,39,39,79,79,79,79,41,41,41,41,79,79,37,37,103,103,75),
(67,67,67,67,67,119,119,32,32,15,15,69,47,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,48,48,48,48,48,48,62,62,26,26,22,22,22,22,22,22,22,22,22,22,22,22,22,22,22,3,61,61,59,59,33,33,39,81,41,41,36,36,36,36,41,41,37,37,123,123,75),
(67,67,67,67,67,119,119,32,32,15,15,47,69,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,48,48,48,48,48,48,62,62,26,26,22,22,22,22,22,22,22,22,22,22,22,22,22,22,3,3,61,3,59,59,33,33,81,81,41,41,36,36,36,36,41,41,37,37,123,123,75),
(67,67,67,67,67,67,67,32,32,42,42,54,54,29,29,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,48,48,62,62,62,62,26,26,35,35,22,22,30,30,23,23,20,23,30,30,20,23,20,23,30,30,60,24,18,18,31,31,39,39,41,41,79,79,79,79,41,41,79,79,37,37,103),
(67,67,67,67,67,67,67,32,32,42,42,54,54,29,29,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,48,48,62,62,62,62,26,26,35,35,22,22,30,30,23,23,23,20,30,30,23,20,23,20,30,30,24,60,18,18,31,45,39,39,41,41,79,79,79,79,41,41,37,79,37,37,103),
(67,67,67,67,67,67,67,119,119,32,32,15,15,69,47,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,48,48,62,62,26,26,35,35,35,35,22,22,30,30,1,1,1,1,1,1,1,1,1,1,1,1,1,1,7,7,25,25,33,33,76,81,37,37,37,37,37,37,41,41,37,37,103),
(67,67,67,67,67,67,67,119,119,32,32,15,15,47,69,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,48,48,62,62,26,26,35,35,35,35,3,3,30,30,1,1,1,1,1,1,1,1,1,1,1,1,1,1,7,7,25,25,33,33,76,81,37,37,37,37,37,37,41,41,37,37,103),
(67,67,67,67,67,67,67,67,67,32,32,42,42,47,47,49,49,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,62,48,26,26,22,22,22,22,3,3,22,22,30,30,20,20,20,20,38,38,20,20,20,20,38,38,20,20,24,24,25,25,33,33,76,81,37,37,123,123,123,123,37,37,123,123,103),
(67,67,67,67,67,67,67,67,67,32,32,42,15,69,54,16,49,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,48,62,26,26,22,22,22,22,22,22,3,3,30,30,20,20,20,20,38,38,20,20,20,20,38,38,20,20,24,24,25,25,33,33,76,39,37,37,123,123,123,123,37,37,123,123,103),
(67,67,67,67,67,67,67,67,67,32,32,42,42,15,15,16,29,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,62,48,26,26,22,22,30,30,7,30,3,22,1,1,1,1,38,38,38,38,1,1,1,1,1,1,1,7,7,7,45,45,51,51,123,123,103,103,75,75,103,103,103,103,103,103,75),
(67,67,67,67,67,67,67,67,67,32,32,42,42,15,59,69,29,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,48,62,26,26,22,22,30,30,30,30,3,3,1,1,1,1,38,38,38,38,38,1,1,1,1,1,7,7,25,25,45,45,51,51,123,123,103,103,75,75,103,103,103,103,103,103,75),
(67,67,67,67,67,67,67,119,119,32,32,15,15,47,47,49,49,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,29,29,22,22,30,30,23,23,22,22,30,30,20,20,20,20,30,30,23,23,23,23,30,30,60,24,18,18,33,33,39,39,123,123,75,75,75,75,75,75,75,75,75,75,75),
(67,67,67,67,67,67,67,119,119,32,32,15,15,47,47,49,49,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,29,29,22,22,30,30,23,23,3,3,30,30,20,20,20,20,30,30,23,20,23,23,30,30,24,60,18,18,33,31,39,39,123,123,75,75,75,75,75,75,75,75,75,75,75),
(67,67,67,67,67,119,119,32,32,15,15,47,47,29,29,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,29,29,22,22,30,30,30,30,22,22,30,30,30,30,30,30,22,3,22,3,22,3,3,3,61,61,59,59,33,33,46,81,37,37,75,75,75,75,75,75,75,75,75,75,75),
(67,67,67,67,67,119,119,32,32,15,42,47,54,29,29,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,29,29,22,22,30,30,30,30,3,3,30,30,30,30,30,30,3,22,3,22,3,22,3,3,61,61,59,59,33,33,46,81,37,37,75,75,75,75,75,75,75,75,75,75,75),
(67,67,67,119,119,32,32,42,15,54,47,29,29,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,29,29,22,22,30,30,7,7,3,3,60,60,60,60,60,60,3,3,7,7,30,7,7,7,25,25,31,33,41,41,36,46,37,37,103,103,75,75,75,75,75,75,75,75,75),
(67,67,67,119,119,32,32,15,42,47,54,29,29,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,29,29,22,22,30,30,30,30,3,3,60,60,60,60,60,60,3,3,30,30,30,30,7,7,25,25,31,31,33,33,36,79,37,37,103,103,75,75,75,75,75,75,75,75,75),
(67,67,67,32,32,42,42,54,54,29,29,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,29,29,22,22,23,60,60,60,3,3,60,60,60,60,60,60,3,3,7,7,23,23,24,24,25,25,31,31,81,46,41,41,37,37,123,123,75,75,75,75,75,75,75,75,75),
(67,67,67,32,32,42,42,54,54,29,29,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,29,29,22,22,23,23,60,60,3,3,60,60,60,60,60,60,3,3,7,30,60,23,24,24,25,25,33,33,81,81,41,41,37,37,123,123,75,75,75,75,75,75,75,75,75),
(67,119,119,32,32,15,15,69,47,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,29,29,22,22,3,3,3,3,3,3,3,3,3,3,3,3,3,3,30,7,7,7,25,7,45,45,51,51,46,46,41,41,79,79,37,37,103,103,103,103,103,103,103,103,75),
(67,119,119,32,32,15,15,47,69,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,29,29,22,22,3,3,3,3,3,3,3,3,3,61,3,61,3,61,7,7,7,7,25,25,45,45,51,51,46,46,41,41,79,79,37,37,103,103,103,103,103,103,103,103,75),
(67,32,32,42,42,54,54,29,29,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,16,16,29,29,29,29,69,47,47,47,47,47,47,47,54,54,30,30,60,60,3,3,60,60,60,60,18,18,31,31,39,39,79,79,79,79,41,41,79,79,37,37,37,37,37,37,123,123,103),
(67,32,32,42,42,54,54,29,29,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,16,16,49,29,29,29,47,69,47,47,47,47,47,47,47,54,30,35,60,60,3,3,60,60,24,60,18,18,31,31,39,39,79,79,79,79,41,41,79,79,37,37,37,37,37,37,123,123,103),
(119,32,32,15,15,69,47,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,16,16,29,29,22,22,22,22,22,22,22,22,22,22,22,22,3,22,3,3,3,3,3,3,3,3,3,61,59,59,31,31,39,39,79,79,37,37,41,41,79,79,79,79,79,79,41,41,37,37,103),
(119,32,32,15,15,47,69,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,16,16,49,29,22,22,22,22,22,22,22,22,22,22,22,22,22,3,3,3,3,3,3,3,3,3,61,3,61,59,31,31,39,39,79,79,37,37,41,41,79,79,79,79,79,79,41,41,37,37,103),
(119,42,42,54,54,29,29,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,20,20,20,20,22,22,30,30,30,30,1,1,1,1,1,1,1,38,1,1,1,30,30,30,30,30,7,7,25,25,45,31,39,51,76,76,37,37,79,79,41,41,41,41,41,41,79,79,37,37,103),
(119,42,32,54,54,29,29,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,20,20,20,20,22,22,30,30,1,30,1,1,1,1,1,1,1,1,1,1,1,1,30,30,30,30,7,7,25,7,31,45,51,39,76,76,37,37,79,79,41,41,41,41,41,41,79,79,37,37,103),
(32,42,42,47,47,49,49,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,16,16,20,20,30,30,3,3,30,30,23,20,20,20,1,1,20,20,20,20,38,38,38,38,20,20,20,20,1,1,24,24,18,18,33,33,39,39,123,123,37,37,79,79,36,36,41,41,79,79,123,123,75),
(32,42,42,47,54,49,49,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,16,16,20,20,30,30,3,3,30,30,20,23,20,20,1,1,20,20,20,20,38,38,38,38,20,20,20,20,1,1,24,24,18,18,33,33,39,76,123,123,37,37,79,79,36,36,41,41,79,79,123,123,75),
(32,42,42,69,47,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,49,49,20,20,30,30,22,3,1,1,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,1,1,7,25,45,45,51,51,123,123,37,37,79,79,41,41,79,79,37,37,103,103,75),
(32,15,42,69,47,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,49,49,20,20,30,30,3,22,1,1,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,1,1,25,25,45,45,51,51,123,123,37,37,79,79,41,41,79,79,37,37,103,103,75),
(32,42,42,47,47,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,29,29,22,22,22,22,22,3,1,1,20,20,20,20,38,38,20,20,20,20,38,38,38,38,20,20,20,20,38,38,20,20,24,20,25,25,33,33,76,81,79,79,79,79,41,41,37,37,123,123,75,75,75),
(32,42,15,47,47,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,29,29,22,22,22,22,3,22,1,1,20,20,20,20,38,38,20,20,20,20,38,38,38,38,20,25,20,20,38,38,20,20,24,24,25,25,33,33,76,76,79,79,36,79,41,41,37,37,123,123,75,75,75),
(32,42,42,47,47,49,49,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,29,29,22,22,30,30,1,30,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,1,1,25,1,25,25,33,33,76,76,36,36,41,41,79,79,37,37,103,103,75,75,75),
(32,42,42,54,54,49,49,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,29,29,22,22,30,30,30,1,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,1,1,7,7,25,25,33,33,76,76,36,36,41,41,79,79,37,37,103,103,75,75,75),
(119,42,42,54,54,29,29,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,29,29,22,22,30,30,20,23,1,1,20,20,20,20,1,1,20,20,20,20,38,38,38,38,20,20,20,20,1,1,23,24,24,18,45,31,51,51,41,41,41,41,41,41,79,79,37,37,75,75,75,75,75),
(119,42,32,54,54,29,29,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,29,29,22,22,30,30,23,20,1,1,20,20,20,20,1,1,20,20,20,20,38,38,38,38,20,20,20,20,1,1,23,20,18,24,45,45,51,51,41,41,41,41,41,41,79,79,37,37,75,75,75,75,75),
(119,32,32,15,15,69,47,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,49,49,22,22,1,30,30,30,1,1,30,30,30,30,30,30,30,30,30,30,1,1,1,1,30,30,30,30,30,30,7,7,25,25,31,33,39,76,36,36,36,36,41,41,79,79,37,37,75,75,75,75,75),
(119,32,32,15,15,47,69,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,49,49,22,22,38,1,30,30,1,1,30,30,30,30,30,30,30,30,30,30,30,1,30,1,30,30,30,30,30,30,7,7,25,25,33,31,39,39,36,36,36,36,41,41,79,79,37,37,75,75,75,75,75),
(67,32,32,42,42,54,54,29,29,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,49,49,22,22,22,22,22,22,22,22,3,3,3,3,3,3,3,3,3,3,22,3,22,3,22,3,3,3,3,3,61,61,45,31,51,51,76,76,36,36,41,41,41,41,36,36,37,37,103,103,75,75,75),
(67,32,32,42,42,54,54,49,29,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,49,49,22,22,22,22,22,22,22,22,3,3,3,3,3,3,3,3,3,3,3,22,3,22,3,22,3,3,3,3,61,61,45,45,51,51,76,76,36,36,41,41,41,41,36,36,37,37,103,103,75,75,75),
(67,119,119,32,32,15,15,47,47,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,49,2,49,16,29,29,69,69,3,3,60,60,3,3,60,60,23,23,23,23,23,23,23,23,23,23,60,24,18,18,31,31,39,39,79,79,79,79,41,41,36,36,41,41,37,37,123,123,75,75,75),
(67,119,119,32,32,15,15,47,69,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,49,49,49,49,29,29,69,69,3,3,60,60,3,3,60,60,23,23,23,23,23,23,23,23,23,23,24,60,18,18,31,31,39,39,79,79,79,79,41,41,36,36,41,41,37,37,123,123,75,75,75),
(67,67,67,32,32,42,42,54,54,69,69,16,16,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,16,16,49,49,29,29,22,22,30,7,3,3,30,30,30,30,1,1,1,1,1,1,1,1,7,7,25,25,31,31,39,39,79,79,41,41,36,36,36,36,41,41,79,79,37,37,123,123,75),
(67,67,67,32,32,42,42,54,54,29,69,16,16,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,16,16,49,49,29,29,22,3,30,7,3,3,30,30,30,30,38,1,1,1,1,1,1,1,7,7,25,25,31,31,39,39,79,79,41,41,36,36,36,36,41,41,79,79,37,37,123,123,75),
(67,67,67,119,119,32,32,42,42,54,54,47,47,49,49,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,49,49,22,22,22,3,3,22,30,30,1,1,20,20,20,20,38,38,20,20,20,20,7,7,45,45,51,51,79,46,41,41,79,79,36,36,36,36,41,41,79,79,37,37,103),
(67,67,67,119,119,32,32,42,42,54,54,69,69,49,49,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,49,49,22,22,22,22,22,3,30,1,1,1,20,20,20,20,38,38,20,20,20,20,25,7,45,45,51,51,46,46,41,41,79,79,36,36,36,36,41,41,79,79,37,37,103),
(67,67,67,67,67,119,119,32,32,42,42,15,15,69,47,49,49,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,29,49,69,69,22,22,1,1,38,38,38,38,38,38,38,38,38,38,38,38,7,7,25,25,31,31,76,81,41,41,36,36,36,36,36,36,41,41,41,41,37,37,103),
(67,67,67,67,67,119,119,32,32,42,42,15,15,69,47,16,49,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,29,29,69,69,22,22,1,1,38,38,38,38,38,38,38,38,38,38,38,38,7,7,25,25,31,31,39,76,41,41,36,36,36,36,36,36,41,41,41,41,37,37,103),
(67,67,67,67,67,67,67,119,119,32,32,42,42,15,15,16,29,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,29,29,22,22,1,1,1,1,20,20,20,20,1,1,20,20,20,20,1,7,24,24,45,31,39,39,41,41,36,36,41,41,41,41,79,79,37,37,123,123,103),
(67,67,67,67,67,67,67,119,119,32,32,42,42,15,15,16,29,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,29,29,22,22,1,1,1,1,20,20,20,20,1,1,20,20,20,20,7,1,18,24,31,45,39,39,41,41,36,36,41,41,41,41,79,79,37,37,123,123,103),
(67,67,67,67,67,67,67,67,67,119,119,32,32,15,15,16,69,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,29,29,22,22,30,30,30,30,1,1,1,1,1,1,1,1,1,1,30,30,7,7,25,25,33,33,46,46,41,41,79,79,79,79,37,37,123,123,103,103,75),
(67,67,67,67,67,67,67,67,67,119,119,32,32,15,15,29,69,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,29,29,22,22,38,1,30,30,38,1,1,1,1,1,1,1,1,1,30,30,7,7,25,25,33,33,81,46,41,41,79,79,79,79,37,37,123,123,103,103,75),
(67,67,67,67,67,67,67,67,67,32,32,42,42,54,47,29,29,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,49,49,22,22,22,22,22,22,22,22,22,22,22,22,22,22,22,22,22,22,22,3,61,61,31,31,39,39,41,41,79,79,37,37,103,103,75,75,75,75,75),
(67,67,67,67,67,67,67,67,67,32,32,42,42,54,54,29,29,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,49,49,22,22,22,22,22,22,22,22,22,22,22,22,22,22,22,22,22,22,3,3,61,61,31,31,39,39,41,41,79,79,37,37,103,103,75,75,75,75,75),
(67,67,67,67,67,67,67,119,119,32,32,15,15,69,69,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,49,16,62,62,26,26,26,26,26,26,26,26,26,26,26,26,26,26,35,35,30,30,59,59,33,33,81,81,37,37,103,103,75,75,75,75,75,75,75),
(67,67,67,67,67,67,67,119,119,32,32,15,15,47,47,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,49,16,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,35,35,30,126,59,59,33,33,81,81,37,37,103,103,75,75,75,75,75,75,75),
(67,67,67,67,67,67,67,119,119,42,42,54,54,29,29,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,62,48,62,62,62,62,62,62,62,62,62,62,62,62,62,62,26,26,1,38,25,25,33,33,76,81,123,123,75,75,75,75,75,75,75,75,75),
(67,67,67,67,67,67,67,119,119,42,32,54,54,29,29,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,48,62,62,62,62,62,62,62,62,62,62,62,62,62,62,62,26,26,126,30,7,7,31,31,81,81,123,123,75,75,75,75,75,75,75,75,75),
(67,67,67,67,67,67,67,32,32,42,42,47,47,49,49,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,16,16,16,16,16,16,16,16,16,16,16,48,48,48,48,26,26,38,38,45,45,51,51,75,75,103,103,75,75,75,75,75,75,75,75,75),
(67,67,67,67,67,67,67,32,32,42,42,47,54,49,49,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,2,16,16,16,16,16,16,16,16,16,16,16,16,48,48,48,48,26,26,38,126,45,45,51,51,75,75,103,103,75,75,75,75,75,75,75,75,75),
(67,67,67,67,67,67,67,32,32,42,42,69,47,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,48,48,48,48,48,48,48,48,48,48,48,48,48,48,48,48,48,48,48,48,26,26,7,1,45,45,39,51,123,103,75,75,75,75,75,75,75,75,75,75,75),
(67,67,67,67,67,67,67,32,32,15,42,69,47,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,48,48,48,48,48,48,48,48,48,48,48,48,48,48,48,48,48,48,62,48,26,26,1,7,45,45,51,39,123,123,75,75,75,75,75,75,75,75,75,75,75),
(67,67,67,67,67,67,67,32,32,42,42,47,47,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,48,48,48,48,48,48,48,48,48,48,48,48,48,48,48,48,48,48,48,48,62,62,38,38,7,7,31,33,76,39,37,37,75,75,75,75,75,75,75,75,75,75,75),
(67,67,67,67,67,67,67,32,32,42,15,47,47,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,48,48,48,48,48,48,48,48,48,48,48,48,48,48,48,48,48,48,48,48,62,62,35,26,7,7,31,31,76,76,37,37,75,75,75,75,75,75,75,75,75,75,75),
(67,67,67,67,67,67,67,32,32,42,42,47,47,49,49,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,48,48,48,48,48,48,62,62,62,62,62,62,62,62,62,62,62,62,62,62,62,62,26,26,1,7,45,45,33,33,76,76,37,37,103,103,75,75,75,75,75,75,75,75,75),
(67,67,67,67,67,67,67,32,32,42,42,54,54,49,49,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,2,48,48,48,48,48,48,62,62,62,62,62,62,62,62,62,62,62,62,62,62,62,62,26,26,30,1,45,45,33,33,76,76,37,37,103,103,75,75,75,75,75,75,75,75,75),
(67,67,67,67,67,67,67,119,119,42,42,54,54,29,29,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,48,48,48,48,62,62,62,62,26,26,26,26,35,35,35,35,35,35,35,35,35,35,30,38,7,7,31,31,39,76,41,41,37,37,123,123,75,75,75,75,75,75,75,75,75),
(67,67,67,67,67,67,67,119,119,42,32,54,54,29,29,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,2,48,48,48,48,62,62,62,62,26,26,26,26,35,35,35,35,35,35,35,35,35,35,35,35,7,7,31,31,39,39,41,41,37,37,123,123,75,75,75,75,75,75,75,75,75),
(67,67,67,67,67,67,67,119,119,32,32,15,15,69,47,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,48,48,48,48,48,48,62,62,26,26,22,22,22,22,22,22,22,22,22,22,22,22,22,3,61,61,45,45,51,51,46,79,41,41,79,79,37,37,103,103,75,75,75,75,75,75,75),
(67,67,67,67,67,67,67,119,119,32,32,15,15,47,69,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,48,48,48,48,48,48,62,62,26,26,22,22,22,22,22,22,22,22,22,22,22,22,3,3,61,61,45,45,51,51,46,46,41,41,79,79,37,37,103,103,75,75,75,75,75,75,75),
(67,67,67,67,67,67,67,67,67,32,32,42,42,54,54,29,29,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,48,48,62,62,62,62,26,26,35,35,22,22,30,30,23,23,20,23,30,30,20,23,23,23,25,25,45,31,39,39,79,79,79,79,41,41,79,79,37,37,103,103,75,75,75,75,75),
(67,67,67,67,67,67,67,67,67,32,32,42,42,54,54,29,29,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,48,48,62,62,62,62,26,26,35,35,22,22,30,30,23,23,23,20,30,30,23,20,23,24,25,25,31,31,39,51,79,79,79,79,41,41,79,79,37,37,103,103,75,75,75,75,75),
(67,67,67,67,67,67,67,67,67,119,119,32,32,15,15,69,47,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,48,48,62,62,26,26,35,35,35,35,22,22,30,30,1,1,1,1,1,1,1,1,7,7,25,7,45,45,51,39,79,79,37,37,41,41,79,79,79,79,37,37,123,123,103,103,75),
(67,67,67,67,67,67,67,67,67,119,119,32,32,15,15,47,69,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,48,48,62,62,26,26,35,35,35,35,3,3,30,30,1,1,1,1,1,1,1,1,7,7,25,25,45,31,39,39,79,79,37,37,41,41,79,79,79,79,37,37,123,123,103,103,75),
(67,67,67,67,67,67,67,67,67,67,67,32,32,42,42,54,54,29,29,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,62,48,26,26,22,22,22,22,3,3,22,22,30,30,20,20,20,20,38,38,20,20,20,20,7,7,45,45,51,51,76,76,37,37,79,79,41,41,41,41,79,79,37,37,123,123,103),
(67,67,67,67,67,67,67,67,67,67,67,32,32,42,42,54,54,69,29,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,48,62,26,26,22,22,22,22,22,22,3,3,30,30,20,20,20,20,38,38,20,20,20,20,25,7,45,45,51,51,76,76,37,37,79,79,41,41,41,41,79,79,37,37,123,123,103),
(67,67,67,67,67,67,67,67,67,67,67,119,119,32,32,42,15,47,54,29,29,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,62,48,26,26,22,22,30,30,7,30,3,22,1,1,1,1,38,38,38,38,1,1,1,1,7,7,25,25,33,33,81,81,37,37,37,37,79,79,36,36,41,41,41,41,37,37,103),
(67,67,67,67,67,67,67,67,67,67,67,119,119,32,32,15,42,54,47,29,29,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,48,62,26,26,22,22,30,30,30,30,3,3,1,1,1,1,38,38,38,38,38,1,1,1,7,7,25,25,33,33,81,81,37,37,37,37,79,79,36,36,41,41,41,41,37,37,103),
(67,67,67,67,67,67,67,67,67,67,67,67,67,119,119,32,32,15,15,54,47,49,49,16,16,2,2,2,2,2,2,2,2,2,2,2,2,16,16,29,29,22,22,30,30,23,23,22,22,30,30,20,20,20,20,30,30,23,23,23,23,7,7,59,59,33,33,81,81,37,37,37,37,37,37,36,36,41,41,79,79,37,37,103),
(67,67,67,67,67,67,67,67,67,67,67,67,67,119,119,32,32,15,15,69,47,16,49,16,16,2,2,2,2,2,2,2,2,2,2,2,2,16,16,29,29,22,22,30,30,23,23,3,3,30,30,20,20,20,20,30,30,23,20,23,23,7,7,59,59,33,33,39,81,79,37,37,37,37,37,36,36,41,41,79,79,37,37,103),
(67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,119,119,42,32,15,15,16,29,16,16,2,2,2,2,2,2,2,2,2,2,2,2,16,16,29,29,22,22,30,30,30,30,22,22,30,30,30,30,30,30,22,3,22,3,3,3,61,61,59,59,33,33,41,41,36,79,79,79,79,79,41,41,79,79,37,37,123,123,75),
(67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,119,119,32,42,15,15,16,29,16,16,2,2,2,2,2,2,2,2,2,2,2,2,16,16,29,29,22,22,30,30,30,30,3,3,30,30,30,30,30,30,3,22,3,22,3,3,61,61,59,59,33,33,41,33,36,79,79,79,79,79,41,41,79,79,37,37,123,123,75),
(67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,119,119,42,42,15,15,16,29,16,16,2,2,2,2,2,2,2,2,2,2,2,2,16,16,29,29,22,22,30,30,7,7,3,3,60,60,60,60,60,60,3,3,7,7,7,7,7,7,20,25,33,33,41,41,36,36,36,36,36,36,41,41,37,37,123,123,75,75,75),
(67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,119,119,32,42,15,15,29,29,16,16,2,2,2,2,2,2,2,2,2,2,2,2,16,16,29,29,22,22,30,30,30,30,3,3,60,60,60,60,60,60,3,3,30,30,7,30,7,7,25,25,33,33,41,41,36,36,36,36,36,36,41,41,37,37,123,123,75,75,75),
(67,67,67,67,67,67,67,67,67,67,67,67,67,119,119,32,32,15,15,47,47,49,49,16,16,2,2,2,2,2,2,2,2,2,2,2,2,16,16,29,29,22,22,23,60,60,60,3,3,60,60,60,60,60,60,3,3,7,7,23,23,18,18,31,31,51,39,46,46,41,41,41,41,41,41,79,79,37,37,103,103,75,75,75),
(67,67,67,67,67,67,67,67,67,67,67,67,67,119,119,32,32,15,42,47,47,49,49,16,16,2,2,2,2,2,2,2,2,2,2,2,2,16,16,29,29,22,22,23,23,60,60,3,3,60,60,60,60,60,60,3,3,7,30,60,23,24,24,45,45,39,39,46,46,41,41,41,41,41,41,79,79,37,37,103,103,75,75,75),
(67,67,67,67,67,67,67,67,67,67,67,67,67,32,32,42,42,54,54,29,29,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,29,29,22,22,3,3,3,3,3,3,3,3,3,3,3,3,3,3,30,7,7,7,25,25,31,31,39,39,79,79,79,79,36,36,41,41,79,79,37,37,75,75,75,75,75),
(67,67,67,67,67,67,67,67,67,67,67,67,67,32,32,42,42,54,54,29,29,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,29,29,22,22,3,3,3,3,3,3,3,3,3,61,3,61,3,61,7,7,7,7,25,25,31,31,39,39,79,79,79,79,36,36,41,41,79,79,37,37,75,75,75,75,75),
(67,67,67,67,67,67,67,67,67,67,67,119,119,32,32,15,15,69,47,16,16,2,2,2,2,2,2,2,2,2,2,2,2,16,16,16,16,29,29,29,29,69,47,47,47,47,47,47,47,54,54,30,30,60,60,3,3,60,60,60,18,18,18,31,31,39,39,37,37,79,79,36,36,41,41,79,79,37,37,75,75,75,75,75),
(67,67,67,67,67,67,67,67,67,67,67,119,119,32,32,15,15,47,69,16,16,2,2,2,2,2,2,2,2,2,2,2,2,16,16,16,16,49,29,29,29,47,69,47,47,47,47,47,47,47,54,30,35,60,60,3,3,60,60,24,60,18,18,31,31,39,39,37,37,79,79,36,36,41,41,79,79,37,37,75,75,75,75,75),
(67,67,67,67,67,67,67,67,67,67,67,32,32,42,42,54,54,29,29,16,16,2,2,2,2,2,2,2,2,2,2,16,16,16,16,29,29,22,22,22,22,22,22,22,22,22,22,22,22,3,22,3,3,3,3,3,3,3,3,3,3,61,61,45,45,39,51,76,76,79,79,41,41,41,41,36,36,37,37,103,103,75,75,75),
(67,67,67,67,67,67,67,67,67,67,67,32,32,42,42,54,54,29,29,16,16,2,2,2,2,2,2,2,2,2,2,16,16,16,16,49,29,22,22,22,22,22,22,22,22,22,22,22,22,22,3,3,3,3,3,3,3,3,3,3,3,61,61,45,31,51,39,76,76,79,79,41,41,41,41,36,36,37,37,103,103,75,75,75),
(67,67,67,67,67,67,67,67,67,119,119,32,32,15,15,69,47,16,16,2,2,2,2,2,2,2,2,2,2,2,2,16,16,20,20,20,20,22,22,30,30,30,30,1,1,1,1,1,1,1,38,1,1,1,30,30,30,30,30,7,7,7,7,25,25,33,31,76,39,36,36,41,41,36,36,41,41,79,79,123,123,75,75,75),
(67,67,67,67,67,67,67,67,67,119,119,32,32,15,15,47,69,16,16,2,2,2,2,2,2,2,2,2,2,2,2,16,16,20,20,20,20,22,22,30,30,1,30,1,1,1,1,1,1,1,1,1,1,1,1,30,30,30,30,30,30,7,7,25,25,31,31,39,81,36,36,41,41,36,36,41,41,79,79,123,123,75,75,75),
(67,67,67,67,67,67,67,67,67,119,119,42,42,54,54,29,29,16,16,2,2,2,2,2,2,2,2,2,2,16,16,16,16,20,20,30,30,3,3,30,30,23,20,20,20,1,1,20,20,20,20,38,38,38,38,20,20,20,20,1,1,23,24,24,18,45,31,51,51,41,41,36,36,41,41,41,41,36,79,37,37,103,103,75),
(67,67,67,67,67,67,67,67,67,119,119,42,32,54,54,29,29,16,16,2,2,2,2,2,2,2,2,2,2,16,16,16,16,20,20,30,30,3,3,30,30,20,23,20,20,1,1,20,20,20,20,38,38,38,38,20,20,20,20,1,1,23,20,24,24,45,45,39,39,41,41,36,36,41,41,41,41,36,79,37,37,103,103,75),
(67,67,67,67,67,67,67,67,67,32,32,42,42,47,47,49,49,2,2,2,2,2,2,2,2,2,2,2,2,16,16,49,49,20,20,30,30,22,3,1,1,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,1,7,7,25,25,31,33,41,41,41,41,36,36,36,36,41,41,37,37,123,123,75),
(67,67,67,67,67,67,67,67,67,32,32,42,42,47,54,49,49,2,2,2,2,2,2,2,2,2,2,2,2,16,16,49,49,20,20,30,30,3,22,1,1,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,7,7,25,25,33,31,41,41,41,41,36,36,36,36,41,41,37,37,123,123,75),
(67,67,67,67,67,67,67,67,67,32,32,42,42,69,47,16,16,2,2,2,2,2,2,2,2,2,2,2,2,16,16,29,29,22,22,22,22,22,3,1,1,20,20,20,20,38,38,20,20,20,20,38,38,38,38,20,20,20,20,38,38,20,20,20,20,25,25,45,31,41,33,41,41,36,36,79,79,41,41,79,79,37,37,103),
(67,67,67,67,67,67,67,67,67,32,32,15,42,69,47,16,16,2,2,2,2,2,2,2,2,2,2,2,2,16,16,29,29,22,22,22,22,3,22,1,1,20,20,20,20,38,38,20,20,20,20,38,38,38,38,20,25,20,20,38,38,20,20,20,20,25,7,45,45,41,33,41,41,36,36,79,79,41,41,37,79,37,37,103),
(67,67,67,67,67,67,67,67,67,32,32,42,42,47,47,16,16,2,2,2,2,2,2,2,2,2,2,2,2,16,16,29,29,22,22,30,30,1,30,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,1,25,7,25,25,41,33,46,46,79,79,37,37,37,37,41,41,37,37,103),
(67,67,67,67,67,67,67,67,67,32,32,42,15,47,47,16,16,2,2,2,2,2,2,2,2,2,2,2,2,16,16,29,29,22,22,30,30,30,1,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,1,38,7,7,25,25,33,33,46,46,79,79,37,37,37,37,41,41,37,37,103),
(67,67,67,67,67,67,67,67,67,32,32,42,42,47,47,49,49,2,2,2,2,2,2,2,2,2,2,2,2,16,16,29,29,22,22,30,30,20,23,1,1,20,20,20,20,1,1,20,20,20,20,38,38,38,38,20,20,20,20,1,1,20,20,20,20,7,7,18,18,41,33,76,81,37,37,123,123,123,123,37,37,123,123,103),
(67,67,67,67,67,67,67,67,67,32,32,42,42,54,54,49,49,2,2,2,2,2,2,2,2,2,2,2,2,16,16,29,29,22,22,30,30,23,20,1,1,20,20,20,20,1,1,20,20,20,20,38,38,38,38,20,20,20,20,1,1,20,20,20,20,7,25,18,18,33,33,76,81,37,37,123,123,123,123,37,37,123,123,103),
(67,67,67,67,67,67,67,67,67,119,119,42,42,54,54,29,29,16,16,2,2,2,2,2,2,2,2,2,2,16,16,49,49,22,22,1,30,30,30,1,1,30,30,30,30,30,30,30,30,30,30,1,1,1,1,30,30,30,30,30,30,30,30,7,7,25,25,45,31,51,51,123,123,103,103,75,75,103,103,103,103,103,103,75),
(67,67,67,67,67,67,67,67,67,119,119,42,32,54,54,29,29,16,16,2,2,2,2,2,2,2,2,2,2,16,16,49,49,22,22,38,1,30,30,1,1,30,30,30,30,30,30,30,30,30,30,30,1,30,1,30,30,30,30,30,30,30,30,7,7,25,7,45,45,51,51,123,123,103,103,75,75,103,103,103,103,103,103,75),
(67,67,67,67,67,67,67,67,67,119,119,32,32,15,15,69,47,16,16,2,2,2,2,2,2,2,2,2,2,16,16,49,49,22,22,22,22,22,22,22,22,3,3,3,3,3,3,3,3,3,3,22,3,22,3,22,3,3,3,3,3,3,3,61,61,59,59,31,33,39,39,123,123,75,75,75,75,75,75,75,75,75,75,75),
(67,67,67,67,67,67,67,67,67,119,119,32,32,15,15,47,69,16,16,2,2,2,2,2,2,2,2,2,2,16,16,49,49,22,22,22,22,22,22,22,22,3,3,3,3,3,3,3,3,3,3,3,22,3,22,3,22,3,3,3,3,3,3,61,3,59,59,33,33,39,39,123,123,75,75,75,75,75,75,75,75,75,75,75),
(67,67,67,67,67,67,67,67,67,67,67,32,32,42,42,54,54,29,29,16,16,2,2,2,2,2,2,2,2,2,2,16,16,49,2,49,16,29,29,69,69,3,3,60,60,3,3,60,60,23,23,23,23,23,23,23,23,23,23,23,23,23,23,24,18,18,18,41,33,81,81,37,37,75,75,75,75,75,75,75,75,75,75,75),
(67,67,67,67,67,67,67,67,67,67,67,32,32,42,42,54,54,29,29,16,16,2,2,2,2,2,2,2,2,2,2,16,16,49,49,49,49,29,29,69,69,3,3,60,60,3,3,60,60,23,23,23,23,23,23,23,23,23,23,23,23,23,23,18,18,18,18,33,33,81,81,37,37,75,75,75,75,75,75,75,75,75,75,75),
(67,67,67,67,67,67,67,67,67,67,67,119,119,32,32,15,15,69,69,16,16,2,2,2,2,2,2,2,2,2,2,2,2,16,16,16,16,49,49,29,29,22,22,30,7,3,3,30,30,30,30,1,1,1,1,1,1,1,1,1,1,7,7,25,25,45,33,33,41,46,46,37,37,103,103,75,75,75,75,75,75,75,75,75),
(67,67,67,67,67,67,67,67,67,67,67,119,119,32,32,15,15,69,69,16,16,2,2,2,2,2,2,2,2,2,2,2,2,16,16,16,16,49,49,29,29,22,3,30,7,3,3,30,30,30,30,38,1,1,1,1,1,1,1,1,1,7,7,25,25,31,31,41,41,46,46,37,37,103,103,75,75,75,75,75,75,75,75,75),
(67,67,67,67,67,67,67,67,67,67,67,67,67,32,32,15,15,47,47,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,49,49,22,22,22,3,3,22,30,30,1,1,20,20,20,20,38,38,20,20,20,20,7,7,25,25,31,31,76,39,41,41,37,37,123,123,75,75,75,75,75,75,75,75,75),
(67,67,67,67,67,67,67,67,67,67,67,67,67,32,32,15,15,69,69,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,49,49,22,22,22,22,22,3,30,1,1,1,20,20,20,20,38,38,20,20,20,20,7,7,25,25,31,33,76,46,41,41,37,37,123,123,75,75,75,75,75,75,75,75,75),
(67,67,67,67,67,67,67,67,67,67,67,119,119,32,32,15,15,29,69,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,29,49,69,69,22,22,1,1,38,38,38,38,38,38,38,38,38,38,1,1,7,25,45,45,51,51,79,46,41,41,79,79,37,37,103,103,103,103,103,103,103,103,75),
(67,67,67,67,67,67,67,67,67,67,67,119,119,32,42,15,15,29,69,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,29,29,69,69,22,22,1,1,38,38,38,38,38,38,38,38,38,38,38,1,7,7,45,45,51,51,79,46,41,41,79,79,37,37,103,103,103,103,103,103,103,103,75),
(67,67,67,67,67,67,67,67,67,119,119,32,32,15,15,47,47,49,49,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,29,29,22,22,1,1,38,38,20,20,20,20,38,38,20,20,20,20,25,25,45,45,51,39,79,79,79,79,41,41,37,37,37,37,123,123,37,37,123,123,103),
(67,67,67,67,67,67,67,67,67,119,119,32,32,42,15,54,54,49,49,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,29,29,22,22,38,1,38,38,20,25,20,20,38,38,20,20,20,20,25,7,45,31,51,51,79,79,79,79,41,41,37,37,37,37,123,123,37,37,123,123,103),
(67,67,67,67,67,67,67,67,67,119,119,42,32,54,54,47,69,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,29,29,22,22,38,38,38,38,38,38,38,38,38,38,38,38,38,1,25,7,45,31,51,76,79,79,79,79,41,41,79,79,37,37,37,37,41,41,37,37,123),
(67,67,67,67,67,67,67,67,67,119,119,32,42,54,54,69,69,16,16,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,16,16,29,29,22,22,38,38,38,38,38,38,38,38,38,38,38,38,38,1,25,25,45,31,39,39,79,79,79,79,41,41,79,79,37,37,37,37,41,41,37,37,123)
);

type pipe_rom is array (0 to PipeWidth, 0 to PipeHeight) of integer range 0 to 127;
constant pipespr : pipe_rom := (
(21,21,21,21,21,21,21,21,21,21,21,21,21,21,21,21,21,21,21,21,21,21,21,21,127,127,127),
(21,21,21,21,21,21,21,21,21,21,21,21,21,21,21,21,21,21,21,21,21,21,21,21,127,127,127),
(21,21,66,66,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,56,56,21,21,21,21,21),
(21,21,66,66,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,56,56,21,21,21,21,21),
(21,21,65,65,68,68,64,64,68,68,64,64,64,64,64,64,64,64,64,64,56,56,21,21,56,56,17),
(21,21,65,65,68,68,64,64,68,68,64,64,64,64,64,64,64,64,64,64,56,56,21,21,56,56,17),
(21,21,12,12,63,63,63,63,63,63,63,63,63,63,63,63,63,63,78,78,56,56,21,21,56,56,8),
(21,21,12,12,63,63,63,63,63,63,63,63,63,63,63,63,63,63,78,78,56,56,21,21,56,56,8),
(21,21,64,64,19,19,19,19,19,19,19,19,19,19,19,19,19,19,19,19,56,56,21,21,56,56,6),
(21,21,64,64,19,19,19,19,19,19,19,19,19,19,19,19,19,19,19,19,56,56,21,21,56,56,6),
(21,21,63,63,63,63,78,78,63,63,63,63,63,63,63,63,78,78,63,63,56,56,21,21,56,56,9),
(21,21,63,63,63,63,78,78,63,63,63,63,63,63,63,63,78,78,63,63,56,56,21,21,56,56,9),
(21,21,19,19,64,64,68,68,64,64,68,68,68,68,64,64,64,64,64,64,56,56,21,21,56,56,13),
(21,21,19,19,64,64,68,68,64,64,68,68,68,68,64,64,64,64,64,64,56,56,21,21,56,56,13),
(21,21,63,63,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,56,56,21,21,56,56,12),
(21,21,63,63,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,56,56,21,21,56,56,12),
(21,21,68,68,65,65,65,65,82,82,82,82,82,82,82,82,65,65,65,65,56,56,21,21,56,56,40),
(21,21,68,68,65,65,65,65,82,82,82,82,82,82,82,82,65,65,65,65,56,56,21,21,56,56,40),
(21,21,12,12,66,66,66,66,66,66,66,66,66,66,66,66,66,66,66,66,56,56,21,21,56,56,19),
(21,21,12,12,66,66,66,66,66,66,66,66,66,66,66,66,66,66,66,66,56,56,21,21,56,56,19),
(21,21,64,64,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,56,56,21,21,56,56,40),
(21,21,64,64,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,56,56,21,21,56,56,40),
(21,21,12,12,124,124,124,124,124,124,124,124,124,124,124,124,124,124,124,124,56,56,21,21,56,56,12),
(21,21,12,12,124,124,124,124,124,124,124,124,124,124,124,124,124,124,124,124,56,56,21,21,56,56,12),
(21,21,65,65,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,56,56,21,21,56,56,13),
(21,21,65,65,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,56,56,21,21,56,56,13),
(21,21,66,66,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,56,56,21,21,56,56,9),
(21,21,66,66,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,56,56,21,21,56,56,9),
(21,21,9,9,74,74,74,74,74,74,74,74,74,74,74,74,74,74,74,74,56,56,21,21,56,56,6),
(21,21,9,9,74,74,74,74,74,74,74,74,74,74,74,74,74,74,74,74,56,56,21,21,56,56,6),
(21,21,124,124,17,17,17,17,17,17,17,17,17,17,17,17,17,17,17,17,56,56,21,21,56,56,8),
(21,21,124,124,17,17,17,17,17,17,17,17,17,17,17,17,17,17,17,17,56,56,21,21,56,56,8),
(21,21,6,6,77,77,77,77,77,77,77,77,77,77,77,77,77,77,77,77,56,56,21,21,56,56,17),
(21,21,6,6,14,77,77,77,77,77,77,77,14,77,77,77,14,77,77,77,56,56,21,21,56,56,17),
(21,21,8,8,14,14,27,14,27,14,27,14,14,14,27,14,14,27,27,14,56,56,21,21,56,56,14),
(21,21,8,8,14,27,14,27,14,27,14,27,14,27,14,27,14,14,14,27,56,56,21,21,56,56,14),
(21,21,74,74,80,27,27,27,80,27,80,27,80,27,80,27,80,80,80,27,56,56,21,21,56,56,27),
(21,21,74,74,80,80,27,27,80,80,80,80,80,80,80,80,80,80,80,80,56,56,21,21,56,56,27),
(21,21,17,17,71,71,71,71,71,71,71,71,71,71,71,71,71,71,71,71,56,56,21,21,56,56,57),
(21,21,17,17,71,71,71,71,71,71,71,71,71,71,71,71,71,71,71,71,56,56,21,21,56,56,57),
(21,21,77,77,70,70,70,70,70,70,70,70,70,70,70,70,70,70,70,70,56,56,21,21,56,56,56),
(21,21,14,77,70,70,70,70,70,70,70,70,70,70,70,70,70,70,70,70,56,56,21,21,56,56,56),
(21,21,14,14,56,56,56,56,56,56,56,56,56,56,56,56,56,56,56,56,56,56,21,21,56,56,56),
(21,21,14,27,56,56,56,56,56,56,56,56,56,56,56,56,56,56,56,56,56,56,21,21,56,56,56),
(21,21,80,80,56,56,56,56,56,56,56,56,56,56,56,56,56,56,56,56,56,56,21,21,56,56,56),
(21,21,80,80,56,56,56,56,56,56,56,56,56,56,56,56,56,56,56,56,56,56,21,21,56,56,56),
(21,21,71,71,56,56,56,56,56,56,56,56,56,56,56,56,56,56,56,56,56,56,21,21,56,56,56),
(21,21,71,71,56,56,56,56,56,56,56,56,56,56,56,56,56,56,56,56,56,56,21,21,56,56,56),
(21,21,70,70,56,56,56,56,56,56,56,56,56,56,56,56,56,56,56,56,56,56,21,21,21,21,21),
(21,21,70,70,56,56,56,56,56,56,56,56,56,56,56,56,56,56,56,56,56,56,21,21,21,21,21),
(21,21,21,21,21,21,21,21,21,21,21,21,21,21,21,21,21,21,21,21,21,21,21,21,127,127,127),
(21,21,21,21,21,21,21,21,21,21,21,21,21,21,21,21,21,21,21,21,21,21,21,21,127,127,127));

type bdp is  array(0 to 1) of std_logic_vector(7 downto 0);

constant BigDigitPalette : bdp := ( x"FF", x"00" );

type bigdigit_rom is array (0 to 9, 0 to BigDigitWidth - 1, 0 to BigDigitHeight - 1) of integer range 0 to 2;
constant bigdigits : bigdigit_rom := (
(
(1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2),
(1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
(1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
(2,2,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
(2,2,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1)),
(
(2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2),
(2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2),
(2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2),
(2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2),
(1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2),
(1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2),
(1,1,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2),
(1,1,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
(1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
(2,2,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
(2,2,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
(2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2),
(2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2),
(2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2),
(2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2)),
(
(1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2),
(1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2),
(1,1,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
(1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
(2,2,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
(2,2,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1)),
(
(1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2),
(1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2),
(1,1,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
(1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
(2,2,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
(2,2,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1)),
(
(1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,2,2,2),
(1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,2,2,2),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,2,2,2,2,2,2),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,2,2,2,2,2,2),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,2,2,2,2,2,2),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,2,2,2,2,2,2),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,2,2,2,2,2,2),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,2,2,2,2,2,2),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,2,2,2,2,2,2),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,2,2,2,2,2,2),
(1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,2,2),
(1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,2,2),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
(1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
(2,2,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
(2,2,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1)),
(
(1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2),
(1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
(1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
(2,2,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
(2,2,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1)),
(
(1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2),
(1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
(1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
(2,2,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
(2,2,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1)),
(
(1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2),
(1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,2,2,2,2,2,2,2,2,2,2,2,2,2,2),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,2,2,2,2,2,2,2,2,2,2,2,2,2,2),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,2,2,2,2,2,2,2,2,2,2,2,2,2,2),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,2,2,2,2,2,2,2,2,2,2,2,2,2,2),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,2,2,2,2,2,2,2,2,2,2,2,2,2,2),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,2,2,2,2,2,2,2,2,2,2,2,2,2,2),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,2,2,2,2,2,2,2,2,2,2,2,2,2,2),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,2,2,2,2,2,2,2,2,2,2,2,2,2,2),
(1,1,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2),
(1,1,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
(1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
(2,2,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
(2,2,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1)),
(
(1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2),
(1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
(1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
(2,2,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
(2,2,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1)),
(
(1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2),
(1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1),
(1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
(1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
(2,2,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
(2,2,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1)));

type bottom_bg_palette_ROM is array (0 to 6) of std_logic_vector(7 downto 0);
constant R_bottom_bg_rom : bottom_bg_palette_ROM := 
	(x"9c",x"73",x"e4",x"55",x"d7",x"54",x"de");

constant G_bottom_bg_rom : bottom_bg_palette_ROM := (
x"e6",x"bf",x"fd",x"80",x"a8",x"38",x"d8");

constant B_bottom_bg_rom : bottom_bg_palette_ROM := (
x"59",
x"2e",
x"8b",
x"22",
x"4c",
x"47",
x"95");


type bottom_bg_rom is array (0 to 23, 0 to 21) of integer range 0 to 6;
constant bottom_bg: bottom_bg_rom := (
(5,4,4,0,0,0,0,0,0,0,0,0,0,0,0,1,1,3,3,2,2,6),
(5,4,4,0,0,0,0,0,0,0,0,0,0,0,0,1,1,3,3,2,2,6),
(5,4,4,0,0,0,0,0,0,0,0,0,0,1,1,1,1,3,3,2,2,6),
(5,4,4,0,0,0,0,0,0,0,0,0,0,1,1,1,1,3,3,2,2,6),
(5,4,4,0,0,0,0,0,0,0,0,1,1,1,1,1,1,3,3,2,2,6),
(5,4,4,0,0,0,0,0,0,0,0,1,1,1,1,1,1,3,3,2,2,6),
(5,4,4,0,0,0,0,0,0,1,1,1,1,1,1,1,1,3,3,2,2,6),
(5,4,4,0,0,0,0,0,0,1,1,1,1,1,1,1,1,3,3,2,2,6),
(5,4,4,0,0,0,0,1,1,1,1,1,1,1,1,1,1,3,3,2,2,6),
(5,4,4,0,0,0,0,1,1,1,1,1,1,1,1,1,1,3,3,2,2,6),
(5,4,4,0,0,1,1,1,1,1,1,1,1,1,1,1,1,3,3,2,2,6),
(5,4,4,0,0,1,1,1,1,1,1,1,1,1,1,1,1,3,3,2,2,6),
(5,4,4,1,1,1,1,1,1,1,1,1,1,1,1,0,0,3,3,2,2,6),
(5,4,4,1,1,1,1,1,1,1,1,1,1,1,1,0,0,3,3,2,2,6),
(5,4,4,1,1,1,1,1,1,1,1,1,1,0,0,0,0,3,3,2,2,6),
(5,4,4,1,1,1,1,1,1,1,1,1,1,0,0,0,0,3,3,2,2,6),
(5,4,4,1,1,1,1,1,1,1,1,0,0,0,0,0,0,3,3,2,2,6),
(5,4,4,1,1,1,1,1,1,1,1,0,0,0,0,0,0,3,3,2,2,6),
(5,4,4,1,1,1,1,1,1,0,0,0,0,0,0,0,0,3,3,2,2,6),
(5,4,4,1,1,1,1,1,1,0,0,0,0,0,0,0,0,3,3,2,2,6),
(5,4,4,1,1,1,1,0,0,0,0,0,0,0,0,0,0,3,3,2,2,6),
(5,4,4,1,1,1,1,0,0,0,0,0,0,0,0,0,0,3,3,2,2,6),
(5,4,4,1,1,0,0,0,0,0,0,0,0,0,0,0,0,3,3,2,2,6),
(5,4,4,1,1,0,0,0,0,0,0,0,0,0,0,0,0,3,3,2,2,6));


type getready_palette_ROM is array (0 to 4) of std_logic_vector(7 downto 0);
constant R_getready_rom : getready_palette_ROM := (
x"ff",x"66", x"66", x"00", x"FF");
constant G_getready_rom : getready_palette_ROM := (
x"ff", x"cc", x"33", x"99", x"FF");
constant B_getready_rom : getready_palette_ROM := (
x"ff", x"66", x"33", x"33", x"FF");

type getready_rom is array (0 to 183, 0 to 49) of integer range 0 to 4;
constant getready: getready_rom := (
(4,4,4,4,4,4,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,4,4,4,4,4,4,4,4,4,4,4,4,4,4),
(4,4,4,4,4,4,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,4,4,4,4,4,4,4,4,4,4,4,4,4,4),
(4,4,4,4,2,2,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,2,2,4,4,4,4,4,4,4,4,4,4,4,4),
(4,4,4,4,2,2,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,2,2,4,4,4,4,4,4,4,4,4,4,4,4),
(4,4,2,2,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,0,0,2,2,4,4,4,4,4,4,4,4,4,4),
(4,4,2,2,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,0,0,2,2,4,4,4,4,4,4,4,4,4,4),
(2,2,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,0,0,2,2,4,4,4,4,4,4,4,4),
(2,2,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,0,0,2,2,4,4,4,4,4,4,4,4),
(2,2,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,2,2,4,4,4,4,4,4,4,4),
(2,2,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,2,2,4,4,4,4,4,4,4,4),
(2,2,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,2,2,4,4,4,4,4,4,4,4),
(2,2,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,2,2,4,4,4,4,4,4,4,4),
(2,2,0,0,1,1,1,1,1,1,3,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,3,3,0,0,2,2,4,4,4,4,4,4,4,4),
(2,2,0,0,1,1,1,1,1,1,3,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,3,3,0,0,2,2,4,4,4,4,4,4,4,4),
(2,2,0,0,1,1,1,1,1,1,3,3,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,2,2,4,4,4,4,4,4,4,4),
(2,2,0,0,1,1,1,1,1,1,3,3,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,2,2,4,4,4,4,4,4,4,4),
(2,2,0,0,1,1,1,1,1,1,3,3,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,2,2,4,4,4,4,4,4,4,4),
(2,2,0,0,1,1,1,1,1,1,3,3,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,2,2,4,4,4,4,4,4,4,4),
(2,2,0,0,1,1,1,1,1,1,3,3,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,2,2,4,4,4,4,4,4,4,4),
(2,2,0,0,1,1,1,1,1,1,3,3,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,2,2,4,4,4,4,4,4,4,4),
(2,2,0,0,1,1,1,1,1,1,3,3,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,2,2,4,4,4,4,4,4,4,4),
(2,2,0,0,1,1,1,1,1,1,3,3,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,2,2,4,4,4,4,4,4,4,4),
(2,2,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,2,2,4,4,4,4,4,4,4,4),
(2,2,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,2,2,4,4,4,4,4,4,4,4),
(2,2,2,2,2,2,2,2,2,2,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,0,0,2,2,2,2,4,4,4,4,4,4,4,4),
(2,2,2,2,2,2,2,2,2,2,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,0,0,2,2,2,2,4,4,4,4,4,4,4,4),
(4,4,4,4,2,2,2,2,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,0,0,2,2,4,4,4,4,4,4,4,4),
(4,4,4,4,2,2,2,2,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,0,0,2,2,4,4,4,4,4,4,4,4),
(4,4,4,4,2,2,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,2,2,4,4,4,4,4,4,4,4),
(4,4,4,4,2,2,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,2,2,4,4,4,4,4,4,4,4),
(4,4,4,4,2,2,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,2,2,4,4,4,4,4,4,4,4),
(4,4,4,4,2,2,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,2,2,4,4,4,4,4,4,4,4),
(4,4,4,4,2,2,0,0,1,1,1,1,1,1,1,1,3,3,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,2,2,4,4,4,4,4,4,4,4),
(4,4,4,4,2,2,0,0,1,1,1,1,1,1,1,1,3,3,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,2,2,4,4,4,4,4,4,4,4),
(4,4,4,4,2,2,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,0,0,0,0,0,0,0,0,2,2,4,4,4,4,4,4,4,4),
(4,4,4,4,2,2,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,0,0,0,0,0,0,0,0,2,2,4,4,4,4,4,4,4,4),
(4,4,4,4,2,2,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,2,2,2,2,2,2,2,2,2,2,4,4,4,4,4,4,4,4),
(4,4,4,4,2,2,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,2,2,2,2,2,2,2,2,2,2,4,4,4,4,4,4,4,4),
(4,4,4,4,4,4,2,2,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,2,2,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4),
(4,4,4,4,4,4,2,2,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,2,2,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4),
(4,4,4,4,4,4,4,4,2,2,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,2,2,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4),
(4,4,4,4,4,4,4,4,2,2,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,2,2,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4),
(4,4,4,4,4,4,4,4,0,0,2,2,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,2,2,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4),
(4,4,4,4,4,4,4,4,0,0,2,2,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,2,2,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4),
(2,2,2,2,2,2,2,2,2,2,2,2,0,0,1,1,1,1,1,1,3,3,0,0,2,2,2,2,2,2,2,2,2,2,2,2,4,4,4,4,4,4,4,4,4,4,4,4,4,4),
(2,2,2,2,2,2,2,2,2,2,2,2,0,0,1,1,1,1,1,1,3,3,0,0,2,2,2,2,2,2,2,2,2,2,2,2,4,4,4,4,4,4,4,4,4,4,4,4,4,4),
(2,2,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,3,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,2,2,4,4,4,4,4,4,4,4,4,4,4,4),
(2,2,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,3,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,2,2,4,4,4,4,4,4,4,4,4,4,4,4),
(2,2,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,0,0,2,2,4,4,4,4,4,4,4,4,4,4),
(2,2,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,0,0,2,2,4,4,4,4,4,4,4,4,4,4),
(2,2,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,0,0,2,2,4,4,4,4,4,4,4,4),
(2,2,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,0,0,2,2,4,4,4,4,4,4,4,4),
(2,2,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,2,2,4,4,4,4,4,4,4,4),
(2,2,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,2,2,4,4,4,4,4,4,4,4),
(2,2,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,2,2,4,4,4,4,4,4,4,4),
(2,2,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,2,2,4,4,4,4,4,4,4,4),
(2,2,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,3,3,0,0,0,0,0,0,0,0,1,1,1,1,1,1,3,3,0,0,2,2,4,4,4,4,4,4,4,4),
(2,2,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,3,3,0,0,0,0,0,0,0,0,1,1,1,1,1,1,3,3,0,0,2,2,4,4,4,4,4,4,4,4),
(2,2,2,2,2,2,2,2,2,2,2,2,0,0,1,1,1,1,1,1,3,3,0,0,2,2,2,2,0,0,1,1,1,1,1,1,3,3,0,0,2,2,4,4,4,4,4,4,4,4),
(2,2,2,2,2,2,2,2,2,2,2,2,0,0,1,1,1,1,1,1,3,3,0,0,2,2,2,2,0,0,1,1,1,1,1,1,3,3,0,0,2,2,4,4,4,4,4,4,4,4),
(4,4,4,4,4,4,4,4,4,4,2,2,0,0,0,0,0,0,0,0,0,0,0,0,2,2,2,2,0,0,0,0,0,0,0,0,0,0,0,0,2,2,4,4,4,4,4,4,4,4),
(4,4,4,4,4,4,4,4,4,4,2,2,0,0,0,0,0,0,0,0,0,0,0,0,2,2,2,2,0,0,0,0,0,0,0,0,0,0,0,0,2,2,4,4,4,4,4,4,4,4),
(4,4,4,4,4,4,4,4,4,4,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,4,4,4,4,4,4,4,4),
(4,4,4,4,4,4,4,4,4,4,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,4,4,4,4,4,4,4,4),
(4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4),
(4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4),
(4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4),
(4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4),
(2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,4,4,4,4,4,4,4,4,4,4),
(2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,4,4,4,4,4,4,4,4,4,4),
(2,2,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,2,2,4,4,4,4,4,4,4,4),
(2,2,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,2,2,4,4,4,4,4,4,4,4),
(2,2,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,2,2,4,4,4,4,4,4,4,4),
(2,2,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,2,2,4,4,4,4,4,4,4,4),
(2,2,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,2,2,4,4,4,4,4,4,4,4),
(2,2,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,2,2,4,4,4,4,4,4,4,4),
(2,2,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,2,2,4,4,4,4,4,4,4,4),
(2,2,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,2,2,4,4,4,4,4,4,4,4),
(2,2,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,2,2,4,4,4,4,4,4,4,4),
(2,2,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,1,1,1,3,3,0,0,2,2,4,4,4,4,4,4,4,4),
(2,2,0,0,1,1,1,1,1,1,3,3,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,2,2,4,4,4,4,4,4,4,4),
(2,2,0,0,1,1,1,1,1,1,3,3,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,2,2,4,4,4,4,4,4,4,4),
(2,2,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,2,2,4,4,4,4,4,4,4,4),
(2,2,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,2,2,4,4,4,4,4,4,4,4),
(2,2,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,2,2,4,4,4,4,4,4,4,4),
(2,2,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,2,2,4,4,4,4,4,4,4,4),
(2,2,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,0,0,1,1,1,1,3,3,0,0,2,2,4,4,4,4,4,4,4,4),
(2,2,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,0,0,1,1,1,1,3,3,0,0,2,2,4,4,4,4,4,4,4,4),
(4,4,2,2,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,0,0,0,0,0,0,1,1,3,3,0,0,2,2,4,4,4,4,4,4,4,4),
(4,4,2,2,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,0,0,0,0,0,0,1,1,3,3,0,0,2,2,4,4,4,4,4,4,4,4),
(4,4,4,4,2,2,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,2,2,4,4,4,4,4,4,4,4),
(4,4,4,4,2,2,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,2,2,4,4,4,4,4,4,4,4),
(4,4,4,4,4,4,2,2,2,2,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,0,0,2,2,2,2,4,4,4,4,4,4,4,4),
(4,4,4,4,4,4,2,2,2,2,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,0,0,2,2,2,2,4,4,4,4,4,4,4,4),
(4,4,4,4,4,4,2,2,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,0,0,2,2,4,4,4,4,4,4,4,4),
(4,4,4,4,4,4,2,2,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,0,0,2,2,4,4,4,4,4,4,4,4),
(4,4,4,4,2,2,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,2,2,4,4,4,4,4,4,4,4),
(4,4,4,4,2,2,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,2,2,4,4,4,4,4,4,4,4),
(4,4,4,4,2,2,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,2,2,4,4,4,4,4,4,4,4),
(4,4,4,4,2,2,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,2,2,4,4,4,4,4,4,4,4),
(4,4,4,4,2,2,0,0,1,1,1,1,1,1,1,1,3,3,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,2,2,4,4,4,4,4,4,4,4),
(4,4,4,4,2,2,0,0,1,1,1,1,1,1,1,1,3,3,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,2,2,4,4,4,4,4,4,4,4),
(4,4,4,4,2,2,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,0,0,0,0,0,0,0,0,2,2,4,4,4,4,4,4,4,4),
(4,4,4,4,2,2,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,0,0,0,0,0,0,0,0,2,2,4,4,4,4,4,4,4,4),
(4,4,4,4,2,2,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,2,2,2,2,2,2,2,2,2,2,4,4,4,4,4,4,4,4),
(4,4,4,4,2,2,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,2,2,2,2,2,2,2,2,2,2,4,4,4,4,4,4,4,4),
(4,4,4,4,4,4,2,2,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,2,2,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4),
(4,4,4,4,4,4,2,2,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,2,2,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4),
(4,4,4,4,4,4,4,4,2,2,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,2,2,2,2,4,4,4,4,4,4,4,4,4,4,4,4,4,4),
(4,4,4,4,4,4,4,4,2,2,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,2,2,2,2,4,4,4,4,4,4,4,4,4,4,4,4,4,4),
(4,4,4,4,4,4,4,4,4,4,2,2,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,2,2,4,4,4,4,4,4,4,4,4,4,4,4),
(4,4,4,4,4,4,4,4,4,4,2,2,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,2,2,4,4,4,4,4,4,4,4,4,4,4,4),
(4,4,4,4,4,4,4,4,4,4,4,4,2,2,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,0,0,2,2,4,4,4,4,4,4,4,4,4,4),
(4,4,4,4,4,4,4,4,4,4,4,4,2,2,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,0,0,2,2,4,4,4,4,4,4,4,4,4,4),
(4,4,4,4,4,4,4,4,4,4,2,2,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,0,0,2,2,4,4,4,4,4,4,4,4),
(4,4,4,4,4,4,4,4,4,4,2,2,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,0,0,2,2,4,4,4,4,4,4,4,4),
(4,4,4,4,4,4,4,4,2,2,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,2,2,4,4,4,4,4,4,4,4),
(4,4,4,4,4,4,4,4,2,2,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,2,2,4,4,4,4,4,4,4,4),
(4,4,4,4,4,4,4,4,2,2,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,2,2,4,4,4,4,4,4,4,4),
(4,4,4,4,4,4,4,4,2,2,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,2,2,4,4,4,4,4,4,4,4),
(4,4,4,4,4,4,4,4,2,2,0,0,1,1,1,1,1,1,1,1,3,3,0,0,0,0,0,0,0,0,1,1,1,1,1,1,3,3,0,0,2,2,4,4,4,4,4,4,4,4),
(4,4,4,4,4,4,4,4,2,2,0,0,1,1,1,1,1,1,1,1,3,3,0,0,0,0,0,0,0,0,1,1,1,1,1,1,3,3,0,0,2,2,4,4,4,4,4,4,4,4),
(4,4,4,4,4,4,4,4,2,2,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,2,2,4,4,4,4,4,4,4,4),
(4,4,4,4,4,4,4,4,2,2,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,2,2,4,4,4,4,4,4,4,4),
(4,4,4,4,4,4,4,4,2,2,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,2,2,4,4,4,4,4,4,4,4),
(4,4,4,4,4,4,4,4,2,2,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,2,2,4,4,4,4,4,4,4,4),
(4,4,4,4,4,4,4,4,2,2,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,2,2,4,4,4,4,4,4,4,4),
(4,4,4,4,4,4,4,4,2,2,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,2,2,4,4,4,4,4,4,4,4),
(4,4,4,4,4,4,4,4,2,2,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,2,2,4,4,4,4,4,4,4,4),
(4,4,4,4,4,4,4,4,2,2,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,2,2,4,4,4,4,4,4,4,4),
(4,4,4,4,4,4,4,4,2,2,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,2,2,4,4,4,4,4,4,4,4),
(4,4,4,4,4,4,4,4,2,2,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,2,2,4,4,4,4,4,4,4,4),
(4,4,4,4,4,4,4,4,2,2,2,2,2,2,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,0,0,2,2,2,2,4,4,4,4,4,4,4,4),
(4,4,4,4,4,4,4,4,2,2,2,2,2,2,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,0,0,2,2,2,2,4,4,4,4,4,4,4,4),
(4,4,4,4,4,4,4,4,4,4,2,2,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,0,0,2,2,4,4,4,4,4,4,4,4),
(4,4,4,4,4,4,4,4,4,4,2,2,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,0,0,2,2,4,4,4,4,4,4,4,4),
(4,4,4,4,4,4,4,4,4,4,2,2,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,2,2,4,4,4,4,4,4,4,4),
(4,4,4,4,4,4,4,4,4,4,2,2,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,2,2,4,4,4,4,4,4,4,4),
(2,2,2,2,2,2,2,2,2,2,2,2,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,2,2,4,4,4,4,4,4,4,4),
(2,2,2,2,2,2,2,2,2,2,2,2,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,2,2,4,4,4,4,4,4,4,4),
(2,2,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,3,3,0,0,0,0,0,0,0,0,1,1,1,1,1,1,3,3,0,0,2,2,4,4,4,4,4,4,4,4),
(2,2,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,3,3,0,0,0,0,0,0,0,0,1,1,1,1,1,1,3,3,0,0,2,2,4,4,4,4,4,4,4,4),
(2,2,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,2,2,4,4,4,4,4,4,4,4),
(2,2,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,2,2,4,4,4,4,4,4,4,4),
(2,2,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,2,2,4,4,4,4,4,4,4,4),
(2,2,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,2,2,4,4,4,4,4,4,4,4),
(2,2,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,2,2,4,4,4,4,4,4,4,4),
(2,2,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,2,2,4,4,4,4,4,4,4,4),
(2,2,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,2,2,4,4,4,4,4,4,4,4),
(2,2,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,2,2,4,4,4,4,4,4,4,4),
(2,2,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,2,2,4,4,4,4,4,4,4,4),
(2,2,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,2,2,4,4,4,4,4,4,4,4),
(2,2,2,2,2,2,2,2,2,2,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,0,0,2,2,2,2,2,2,2,2,4,4,4,4,4,4,4,4),
(2,2,2,2,2,2,2,2,2,2,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,0,0,2,2,2,2,2,2,2,2,4,4,4,4,4,4,4,4),
(4,4,4,4,4,4,4,4,2,2,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,0,0,2,2,2,2,2,2,2,2,2,2,2,2,2,2),
(4,4,4,4,4,4,4,4,2,2,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,0,0,2,2,2,2,2,2,2,2,2,2,2,2,2,2),
(4,4,4,4,4,4,4,4,2,2,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,2,2),
(4,4,4,4,4,4,4,4,2,2,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,2,2),
(4,4,4,4,4,4,4,4,2,2,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,0,0,1,1,1,1,1,1,3,3,0,0,2,2),
(4,4,4,4,4,4,4,4,2,2,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,0,0,1,1,1,1,1,1,3,3,0,0,2,2),
(4,4,4,4,4,4,4,4,2,2,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,3,3,0,0,0,0,1,1,1,1,1,1,3,3,0,0,2,2),
(4,4,4,4,4,4,4,4,2,2,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,3,3,0,0,0,0,1,1,1,1,1,1,3,3,0,0,2,2),
(4,4,4,4,4,4,4,4,2,2,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,2,2),
(4,4,4,4,4,4,4,4,2,2,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,2,2),
(4,4,4,4,4,4,4,4,2,2,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,2,2),
(4,4,4,4,4,4,4,4,2,2,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,2,2),
(4,4,4,4,4,4,4,4,2,2,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,0,0,2,2),
(4,4,4,4,4,4,4,4,2,2,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,0,0,2,2),
(2,2,2,2,2,2,2,2,2,2,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,0,0,2,2,4,4),
(2,2,2,2,2,2,2,2,2,2,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,0,0,2,2,4,4),
(2,2,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,2,2,4,4,4,4),
(2,2,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,2,2,4,4,4,4),
(2,2,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,0,0,1,1,1,1,1,1,3,3,0,0,2,2,2,2,4,4,4,4,4,4),
(2,2,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,0,0,1,1,1,1,1,1,3,3,0,0,2,2,2,2,4,4,4,4,4,4),
(2,2,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,0,0,1,1,1,1,1,1,3,3,0,0,2,2,4,4,4,4,4,4,4,4),
(2,2,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,0,0,1,1,1,1,1,1,3,3,0,0,2,2,4,4,4,4,4,4,4,4),
(2,2,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,0,0,1,1,1,1,1,1,3,3,0,0,2,2,4,4,4,4,4,4,4,4),
(2,2,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,0,0,1,1,1,1,1,1,3,3,0,0,2,2,4,4,4,4,4,4,4,4),
(2,2,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,0,0,1,1,1,1,1,1,3,3,0,0,2,2,4,4,4,4,4,4,4,4),
(2,2,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,3,3,0,0,0,0,1,1,1,1,1,1,3,3,0,0,2,2,4,4,4,4,4,4,4,4),
(2,2,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,2,2,4,4,4,4,4,4,4,4),
(2,2,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,2,2,4,4,4,4,4,4,4,4),
(2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,4,4,4,4,4,4,4,4),
(2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,4,4,4,4,4,4,4,4));

type gameover_palette_ROM is array (0 to 4) of std_logic_vector(7 downto 0);
constant R_gameover_rom : gameover_palette_ROM := (
x"fc",x"ff", x"54", x"e4", x"ff");
constant G_gameover_rom : gameover_palette_ROM := (
x"a0",
x"ff",
x"38",
x"60",
x"ff");
constant B_gameover_rom : gameover_palette_ROM := (
x"48",
x"ff",
x"47",
x"18",
x"ff");

type gameover_rom is array (0 to 191, 0 to 41) of integer range 0 to 4;
constant gameover: gameover_rom := (
(4,4,4,4,4,4,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,4,4,4,4,4,4),
(4,4,4,4,4,4,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,4,4,4,4,4,4),
(4,4,4,4,2,2,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,4,4,4,4),
(4,4,4,4,2,2,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,4,4,4,4),
(4,4,2,2,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,1,1,2,2,4,4),
(4,4,2,2,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,1,1,2,2,4,4),
(2,2,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,1,1,2,2),
(2,2,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,1,1,2,2),
(2,2,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,2,2),
(2,2,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,2,2),
(2,2,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,2,2),
(2,2,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,2,2),
(2,2,1,1,0,0,0,0,0,0,3,3,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,3,3,1,1,2,2),
(2,2,1,1,0,0,0,0,0,0,3,3,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,3,3,1,1,2,2),
(2,2,1,1,0,0,0,0,0,0,3,3,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,2,2),
(2,2,1,1,0,0,0,0,0,0,3,3,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,2,2),
(2,2,1,1,0,0,0,0,0,0,3,3,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,2,2),
(2,2,1,1,0,0,0,0,0,0,3,3,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,2,2),
(2,2,1,1,0,0,0,0,0,0,3,3,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,2,2),
(2,2,1,1,0,0,0,0,0,0,3,3,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,2,2),
(2,2,1,1,0,0,0,0,0,0,3,3,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,2,2),
(2,2,1,1,0,0,0,0,0,0,3,3,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,2,2),
(2,2,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2),
(2,2,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2),
(2,2,2,2,2,2,2,2,2,2,2,2,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,1,1,2,2,2,2),
(2,2,2,2,2,2,2,2,2,2,2,2,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,1,1,2,2,2,2),
(4,4,4,4,4,4,4,4,2,2,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,1,1,2,2),
(4,4,4,4,4,4,4,4,2,2,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,1,1,2,2),
(4,4,4,4,4,4,4,4,2,2,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,2,2),
(4,4,4,4,4,4,4,4,2,2,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,2,2),
(4,4,4,4,4,4,4,4,2,2,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,2,2),
(4,4,4,4,4,4,4,4,2,2,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,2,2),
(4,4,4,4,4,4,4,4,2,2,1,1,0,0,0,0,0,0,0,0,3,3,1,1,1,1,1,1,1,1,0,0,0,0,0,0,3,3,1,1,2,2),
(4,4,4,4,4,4,4,4,2,2,1,1,0,0,0,0,0,0,0,0,3,3,1,1,1,1,1,1,1,1,0,0,0,0,0,0,3,3,1,1,2,2),
(4,4,4,4,4,4,4,4,2,2,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,2,2),
(4,4,4,4,4,4,4,4,2,2,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,2,2),
(4,4,4,4,4,4,4,4,2,2,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,2,2),
(4,4,4,4,4,4,4,4,2,2,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,2,2),
(4,4,4,4,4,4,4,4,2,2,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,2,2),
(4,4,4,4,4,4,4,4,2,2,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,2,2),
(4,4,4,4,4,4,4,4,2,2,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,2,2),
(4,4,4,4,4,4,4,4,2,2,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,2,2),
(4,4,4,4,4,4,4,4,2,2,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2),
(4,4,4,4,4,4,4,4,2,2,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2),
(4,4,4,4,4,4,4,4,2,2,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,2,2),
(4,4,4,4,4,4,4,4,2,2,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,2,2),
(4,4,4,4,4,4,4,4,2,2,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,2,2),
(4,4,4,4,4,4,4,4,2,2,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,2,2),
(4,4,4,4,4,4,4,4,2,2,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,2,2),
(4,4,4,4,4,4,4,4,2,2,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,2,2),
(4,4,4,4,4,4,4,4,2,2,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,2,2),
(4,4,4,4,4,4,4,4,2,2,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,2,2),
(4,4,4,4,4,4,4,4,2,2,1,1,0,0,0,0,0,0,0,0,3,3,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2),
(4,4,4,4,4,4,4,4,2,2,1,1,0,0,0,0,0,0,0,0,3,3,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2),
(4,4,4,4,4,4,4,4,2,2,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,2,2),
(4,4,4,4,4,4,4,4,2,2,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,2,2),
(4,4,4,4,4,4,4,4,2,2,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,2,2),
(4,4,4,4,4,4,4,4,2,2,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,2,2),
(4,4,4,4,4,4,4,4,2,2,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,2,2),
(4,4,4,4,4,4,4,4,2,2,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,2,2),
(4,4,4,4,4,4,4,4,2,2,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,2,2),
(4,4,4,4,4,4,4,4,2,2,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,2,2),
(4,4,4,4,4,4,4,4,2,2,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,2,2),
(4,4,4,4,4,4,4,4,2,2,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,2,2),
(4,4,4,4,4,4,4,4,2,2,1,1,0,0,0,0,0,0,0,0,3,3,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2),
(4,4,4,4,4,4,4,4,2,2,1,1,0,0,0,0,0,0,0,0,3,3,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2),
(4,4,4,4,4,4,4,4,2,2,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,2,2),
(4,4,4,4,4,4,4,4,2,2,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,2,2),
(4,4,4,4,4,4,4,4,2,2,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,2,2),
(4,4,4,4,4,4,4,4,2,2,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,2,2),
(4,4,4,4,4,4,4,4,2,2,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,2,2),
(4,4,4,4,4,4,4,4,2,2,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,2,2),
(4,4,4,4,4,4,4,4,2,2,2,2,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,2,2),
(4,4,4,4,4,4,4,4,2,2,2,2,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,2,2),
(4,4,4,4,4,4,4,4,2,2,2,2,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2),
(4,4,4,4,4,4,4,4,2,2,2,2,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2),
(4,4,4,4,4,4,2,2,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,1,1,2,2,2,2),
(4,4,4,4,4,4,2,2,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,1,1,2,2,2,2),
(4,4,4,4,2,2,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,1,1,2,2),
(4,4,4,4,2,2,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,1,1,2,2),
(4,4,4,4,2,2,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,2,2),
(4,4,4,4,2,2,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,2,2),
(4,4,4,4,2,2,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,2,2),
(4,4,4,4,2,2,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,2,2),
(4,4,4,4,2,2,1,1,0,0,0,0,0,0,0,0,0,0,1,1,1,1,3,3,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,2,2),
(4,4,4,4,2,2,1,1,0,0,0,0,0,0,0,0,0,0,1,1,1,1,3,3,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,2,2),
(4,4,4,4,2,2,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,1,1,1,1,1,1,1,1,2,2),
(4,4,4,4,2,2,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,1,1,1,1,1,1,1,1,2,2),
(4,4,4,4,2,2,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,2,2,2,2,2,2,2,2,2,2),
(4,4,4,4,2,2,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,2,2,2,2,2,2,2,2,2,2),
(4,4,4,4,2,2,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,2,2,4,4,4,4,4,4,4,4),
(4,4,4,4,2,2,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,2,2,4,4,4,4,4,4,4,4),
(4,4,4,4,4,4,2,2,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,2,2,4,4,4,4,4,4,4,4),
(4,4,4,4,4,4,2,2,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,2,2,4,4,4,4,4,4,4,4),
(4,4,4,4,4,4,4,4,2,2,2,2,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,4,4,4,4,4,4,4,4),
(4,4,4,4,4,4,4,4,2,2,2,2,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,4,4,4,4,4,4,4,4),
(4,4,4,4,4,4,4,4,4,4,4,4,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,4,4,4,4,4,4,4,4),
(4,4,4,4,4,4,4,4,4,4,4,4,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,4,4,4,4,4,4,4,4),
(4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4),
(4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4),
(4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4),
(4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4),
(4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4),
(4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4),
(4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4),
(4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4),
(4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4),
(4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4),
(4,4,4,4,4,4,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,4,4,4,4,4,4),
(4,4,4,4,4,4,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,4,4,4,4,4,4),
(4,4,4,4,2,2,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,4,4,4,4),
(4,4,4,4,2,2,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,4,4,4,4),
(4,4,2,2,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,1,1,2,2,4,4),
(4,4,2,2,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,1,1,2,2,4,4),
(2,2,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,1,1,2,2),
(2,2,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,1,1,2,2),
(2,2,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,2,2),
(2,2,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,2,2),
(2,2,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,2,2),
(2,2,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,2,2),
(2,2,1,1,0,0,0,0,0,0,3,3,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,3,3,1,1,2,2),
(2,2,1,1,0,0,0,0,0,0,3,3,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,3,3,1,1,2,2),
(2,2,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,2,2),
(2,2,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,2,2),
(2,2,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,2,2),
(2,2,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,2,2),
(2,2,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,1,1,2,2),
(2,2,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,1,1,2,2),
(4,4,2,2,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,1,1,2,2,2,2),
(4,4,2,2,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,1,1,2,2,2,2),
(4,4,4,4,2,2,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2),
(4,4,4,4,2,2,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2),
(4,4,4,4,4,4,2,2,2,2,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,2,2),
(4,4,4,4,4,4,2,2,2,2,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,2,2),
(4,4,4,4,4,4,4,4,2,2,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,2,2),
(4,4,4,4,4,4,4,4,2,2,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,2,2),
(4,4,4,4,4,4,4,4,2,2,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,2,2),
(4,4,4,4,4,4,4,4,2,2,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,2,2),
(4,4,4,4,4,4,4,4,2,2,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,2,2),
(4,4,4,4,4,4,4,4,2,2,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,2,2),
(4,4,4,4,4,4,4,4,2,2,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,3,3,1,1,2,2),
(4,4,4,4,4,4,4,4,2,2,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,3,3,1,1,2,2),
(4,4,4,4,4,4,4,4,2,2,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,1,1,2,2),
(4,4,4,4,4,4,4,4,2,2,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,1,1,2,2),
(4,4,4,4,4,4,4,4,2,2,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,1,1,2,2,4,4),
(4,4,4,4,4,4,4,4,2,2,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,1,1,2,2,4,4),
(4,4,4,4,4,4,4,4,2,2,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,1,1,2,2,4,4,4,4),
(4,4,4,4,4,4,4,4,2,2,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,1,1,2,2,4,4,4,4),
(4,4,4,4,4,4,4,4,2,2,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,1,1,2,2,4,4,4,4,4,4),
(4,4,4,4,4,4,4,4,2,2,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,1,1,2,2,4,4,4,4,4,4),
(4,4,4,4,4,4,4,4,2,2,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,4,4,4,4),
(4,4,4,4,4,4,4,4,2,2,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,4,4,4,4),
(4,4,4,4,4,4,2,2,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,1,1,2,2,4,4),
(4,4,4,4,4,4,2,2,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,1,1,2,2,4,4),
(4,4,4,4,2,2,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,1,1,2,2),
(4,4,4,4,2,2,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,1,1,2,2),
(4,4,4,4,2,2,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,2,2),
(4,4,4,4,2,2,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,2,2),
(4,4,4,4,2,2,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,2,2),
(4,4,4,4,2,2,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,2,2),
(4,4,4,4,2,2,1,1,0,0,0,0,0,0,0,0,3,3,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,2,2),
(4,4,4,4,2,2,1,1,0,0,0,0,0,0,0,0,3,3,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,2,2),
(4,4,4,4,2,2,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,1,1,1,1,1,1,1,1,2,2),
(4,4,4,4,2,2,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,1,1,1,1,1,1,1,1,2,2),
(4,4,4,4,2,2,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,2,2,2,2,2,2,2,2,2,2),
(4,4,4,4,2,2,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,2,2,2,2,2,2,2,2,2,2),
(4,4,4,4,2,2,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,2,2,4,4,4,4,4,4,4,4),
(4,4,4,4,2,2,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,2,2,4,4,4,4,4,4,4,4),
(4,4,4,4,4,4,2,2,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,2,2,2,2,2,2,2,2,2,2),
(4,4,4,4,4,4,2,2,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,2,2,2,2,2,2,2,2,2,2),
(4,4,4,4,4,4,4,4,2,2,2,2,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2),
(4,4,4,4,4,4,4,4,2,2,2,2,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2),
(4,4,4,4,4,4,4,4,4,4,2,2,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,2,2),
(4,4,4,4,4,4,4,4,4,4,2,2,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,2,2),
(4,4,4,4,4,4,4,4,2,2,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,2,2),
(4,4,4,4,4,4,4,4,2,2,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,2,2),
(4,4,4,4,4,4,4,4,2,2,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,2,2),
(4,4,4,4,4,4,4,4,2,2,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,2,2),
(4,4,4,4,4,4,4,4,2,2,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,2,2),
(4,4,4,4,4,4,4,4,2,2,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,1,1,2,2),
(4,4,4,4,4,4,4,4,2,2,1,1,0,0,0,0,0,0,0,0,3,3,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2),
(4,4,4,4,4,4,4,4,2,2,1,1,0,0,0,0,0,0,0,0,3,3,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2),
(4,4,4,4,4,4,4,4,2,2,1,1,0,0,0,0,0,0,0,0,3,3,1,1,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2),
(4,4,4,4,4,4,4,4,2,2,1,1,0,0,0,0,0,0,0,0,3,3,1,1,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2),
(4,4,4,4,4,4,4,4,2,2,1,1,0,0,0,0,0,0,0,0,3,3,1,1,2,2,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4),
(4,4,4,4,4,4,4,4,2,2,1,1,0,0,0,0,0,0,0,0,3,3,1,1,2,2,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4),
(4,4,4,4,4,4,4,4,2,2,1,1,0,0,0,0,0,0,0,0,3,3,1,1,2,2,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4),
(4,4,4,4,4,4,4,4,2,2,1,1,0,0,0,0,0,0,0,0,3,3,1,1,2,2,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4),
(4,4,4,4,4,4,4,4,2,2,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4),
(4,4,4,4,4,4,4,4,2,2,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4),
(4,4,4,4,4,4,4,4,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4),
(4,4,4,4,4,4,4,4,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4));

type bg16col_palette_ROM is array (0 to 15) of std_logic_vector(7 downto 0);
constant R_bg16col_rom : bg16col_palette_ROM := (
x"d2",
x"e9",
x"9b",
x"cd",
x"ab",
x"a1",
x"b5",
x"62",
x"d5",
x"52",
x"5d",
x"da",
x"e3",
x"df",
x"5e",
x"4f");
constant G_bg16col_rom : bg16col_palette_ROM := (
x"ef",
x"fc",
x"da",
x"ec",
x"e3",
x"dc",
x"e5",
x"cc",
x"f0",
x"cb",
x"c7",
x"f7",
x"fa",
x"f0",
x"df",
x"c1");
constant B_bg16col_rom : bg16col_palette_ROM := (
x"c6",x"d9",
x"d5",x"c4",
x"ba",x"d7",
x"c4",x"7c",
x"c6",x"6c",
x"cc",x"d8",
x"d8",x"cf",
x"70",x"ca");

type bg16col_rom is array (0 to 287, 0 to 83) of integer range 0 to 15;
constant bg16col: bg16col_rom := (
(15,15,15,15,15,15,15,15,15,15,15,10,10,10,10,1,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,1,12,12,5,5,6,6,2,2,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,2,2,2,2,2,2,7,9,14,14,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,10,10,10,1,12,1,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,12,12,5,2,6,6,2,2,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,2,2,2,2,2,2,9,7,14,14,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,10,10,1,11,1,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,1,12,12,5,5,3,3,2,2,0,3,0,0,8,0,8,0,8,0,8,0,8,0,8,0,0,3,3,3,6,3,9,7,14,14,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,10,10,12,11,12,12,1,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,12,12,5,5,3,0,2,2,3,0,0,0,8,8,0,8,0,0,0,8,0,8,0,0,3,0,3,3,3,6,7,7,14,14,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,10,10,11,11,12,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,1,12,12,5,5,5,2,2,2,0,0,0,0,6,6,6,6,8,8,6,6,6,6,8,0,5,5,2,2,3,3,7,7,14,14,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,10,10,11,11,11,12,1,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,12,12,5,5,5,5,5,5,3,0,0,0,6,6,6,6,8,8,6,6,6,6,8,0,5,5,2,5,3,3,7,7,14,14,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,10,10,10,12,11,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,1,12,12,11,12,5,5,0,0,8,8,8,8,8,8,8,8,8,8,8,8,8,8,0,0,3,3,3,6,3,6,9,7,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,10,10,12,11,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,12,12,12,11,5,5,0,0,8,8,8,8,8,8,8,8,8,8,8,8,8,8,0,0,0,3,3,3,3,3,9,7,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,10,10,11,11,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,1,12,12,5,5,0,0,0,0,6,6,6,6,8,0,6,6,6,6,8,0,2,5,2,2,3,6,7,7,9,9,14,14,14,14,14,14,9,9,14,14,14),
(15,15,15,15,15,15,10,10,10,11,11,12,12,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,12,12,5,5,0,0,0,0,6,6,6,6,8,0,6,6,6,6,8,0,5,2,2,2,3,3,7,7,9,7,14,14,14,14,14,14,9,9,14,14,14),
(15,15,15,15,15,15,15,10,10,12,11,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,1,12,12,5,5,0,0,0,3,8,0,8,0,8,0,8,0,8,0,0,3,3,3,3,3,7,7,14,14,14,14,9,9,14,14,9,9,14,14,14,14,14),
(15,15,15,15,15,15,15,10,10,12,11,1,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,12,12,5,5,8,0,3,0,8,0,0,0,0,0,0,0,0,0,3,0,3,3,3,4,7,7,14,14,14,14,9,9,14,14,9,9,14,14,14,14,14),
(15,15,15,15,15,10,10,11,11,12,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,1,12,12,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,2,2,2,2,9,7,14,14,14,14,9,9,14,14,9,9,14,14,14,14,14),
(15,15,15,15,15,10,15,11,11,11,12,1,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,12,12,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,2,5,2,2,2,2,9,7,14,14,14,14,9,9,14,14,9,9,14,14,14,14,14),
(15,15,15,15,15,10,10,11,11,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,1,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,8,13,0,3,0,7,7,14,14,14,14,14,14,14,14,9,9,14,14,14,14,14,14,14),
(15,15,15,15,15,10,10,11,11,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,3,3,7,7,14,14,14,14,14,14,14,14,9,9,14,14,14,14,14,14,14),
(15,15,15,15,10,10,10,12,11,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,1,13,13,13,13,13,13,13,13,13,13,13,13,13,13,0,0,3,3,7,7,14,14,14,14,14,14,14,14,9,9,14,14,14,14,14,14,14),
(15,15,15,15,15,10,10,11,11,1,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,3,0,7,7,14,14,14,14,14,14,14,14,9,9,14,14,14,14,14,14,14),
(15,15,15,15,15,10,10,11,11,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,13,13,13,13,13,13,13,13,13,13,13,13,13,13,0,0,7,7,14,14,14,14,14,14,14,14,9,9,14,14,14,14,14,14,14,14,14),
(15,15,15,15,10,10,10,11,11,1,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,1,13,13,13,13,13,13,13,13,13,13,13,13,13,13,8,0,7,7,14,14,14,14,14,14,14,14,9,9,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,10,10,11,11,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,1,12,1,12,1,12,1,12,1,12,13,13,0,0,7,7,14,14,14,14,14,14,14,14,9,9,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,10,10,11,11,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,1,12,1,1,1,1,1,1,1,1,1,1,1,13,13,0,3,7,7,14,14,14,14,14,14,14,14,9,9,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,10,10,11,11,11,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,0,0,7,7,14,14,14,14,14,14,14,14,9,9,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,10,15,11,12,12,12,1,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,0,3,7,7,14,14,14,14,14,14,14,14,9,9,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,10,10,12,11,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,8,8,7,7,14,14,14,14,14,14,14,14,9,9,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,10,10,10,12,11,1,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,8,3,7,7,14,14,14,14,14,14,14,14,9,9,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,10,10,11,11,11,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,8,13,3,0,7,7,14,14,14,14,14,14,14,14,9,9,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,10,10,11,12,12,12,1,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,1,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,3,3,3,7,7,14,14,14,14,14,14,14,14,9,9,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,10,10,12,11,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,13,13,13,13,13,13,13,13,13,13,13,13,13,13,8,13,13,0,13,13,0,0,13,3,3,3,7,7,14,14,14,14,14,14,9,9,9,9,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,10,10,10,12,11,1,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,1,13,13,13,13,13,13,13,13,13,13,13,13,0,13,13,8,13,13,0,13,13,13,3,13,3,3,7,7,14,14,14,14,14,14,9,9,9,9,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,10,10,11,11,12,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,13,13,13,13,13,13,13,13,13,13,5,5,5,5,5,5,2,5,2,5,5,5,2,5,5,2,2,2,2,2,9,9,9,9,9,9,14,14,14,14,9,9,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,10,10,11,11,12,11,1,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,13,13,13,13,13,13,13,13,13,13,2,5,5,5,5,5,5,5,5,5,5,5,5,5,2,5,2,2,2,10,7,7,9,7,9,9,14,14,14,14,9,9,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,10,10,11,11,12,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,13,13,13,13,13,13,13,13,8,13,5,5,0,0,6,6,6,6,0,3,6,6,6,6,0,3,2,2,2,2,7,9,7,9,9,9,14,14,14,14,9,9,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,10,10,11,12,12,12,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,13,13,13,13,13,13,13,13,13,3,5,5,3,3,6,6,6,6,3,0,6,6,6,6,3,3,2,2,2,2,9,7,9,9,9,9,14,14,14,14,9,9,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,10,15,10,10,11,11,12,12,12,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,13,13,13,13,13,13,8,0,13,13,5,5,0,0,0,0,0,0,8,0,0,0,0,8,0,0,3,3,3,3,3,4,7,7,14,14,14,14,14,14,14,14,9,9,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,15,10,10,12,12,11,11,1,1,1,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,13,13,13,13,13,13,13,13,0,13,2,2,3,0,0,8,0,8,0,0,0,8,0,8,0,0,0,0,3,6,4,3,9,9,14,14,14,14,14,14,14,14,9,9,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,15,10,15,10,10,11,11,11,11,12,12,12,12,12,12,1,1,1,1,1,1,1,1,1,1,13,13,13,13,5,5,2,5,2,2,5,5,0,3,6,6,6,6,8,8,6,6,6,6,8,0,2,2,2,2,3,3,9,7,14,14,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,10,10,11,11,11,1,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,13,13,13,13,5,5,5,5,5,5,2,2,3,0,6,6,6,6,8,8,6,6,6,6,8,0,5,5,2,2,6,3,9,7,14,14,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,10,15,10,10,10,10,11,11,11,11,12,12,1,1,1,1,1,1,1,1,1,1,13,13,13,13,5,5,0,0,3,3,2,5,0,0,8,0,8,8,8,8,8,0,8,0,0,0,3,3,3,3,7,7,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,10,10,10,10,12,11,12,11,12,1,12,12,1,1,1,1,1,1,1,1,13,13,13,13,5,5,3,3,0,0,2,2,0,0,0,8,8,8,8,8,8,0,0,0,0,0,3,3,6,8,7,7,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,10,15,10,10,10,2,11,12,1,1,1,1,1,1,1,1,1,1,1,1,12,12,5,5,0,0,6,6,5,5,0,0,6,6,6,6,0,3,6,6,6,6,3,3,2,2,2,10,7,7,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,10,10,10,10,12,12,12,12,1,1,1,1,1,1,1,1,12,12,12,12,5,5,3,0,6,6,2,2,3,3,6,6,6,6,0,0,6,6,6,6,3,0,2,2,2,4,9,7,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,10,10,1,12,1,1,1,1,1,1,1,1,1,1,1,1,12,12,5,5,0,3,0,0,5,5,0,0,0,0,8,0,5,2,5,2,2,2,2,2,2,2,2,10,7,9,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,10,2,11,11,12,12,1,1,1,1,1,1,1,1,12,12,12,12,5,5,3,0,3,0,2,2,3,3,0,3,0,3,2,5,2,5,2,2,2,2,2,2,2,2,9,7,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,10,10,10,11,12,1,1,1,1,1,1,1,1,1,1,1,1,12,12,5,5,0,0,3,3,2,2,6,6,6,6,6,6,2,2,3,3,0,3,3,3,3,6,9,7,9,9,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,10,10,1,11,12,12,1,1,1,1,1,1,1,1,12,12,12,12,5,5,3,3,0,3,2,2,6,4,6,6,6,6,2,2,0,0,3,0,3,0,3,3,7,7,7,9,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,10,10,11,11,12,12,1,1,1,1,1,1,1,1,1,1,1,1,12,12,5,5,6,6,6,6,2,2,6,6,6,6,4,6,2,2,3,3,6,6,4,4,3,6,7,7,14,14,9,9,14,14,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,10,10,10,11,11,11,12,12,12,1,1,1,1,1,1,1,1,12,12,12,12,5,5,6,6,6,6,2,2,6,6,4,6,6,6,2,2,3,0,6,6,6,4,3,3,9,7,14,14,9,9,14,14,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,10,10,12,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,12,12,5,5,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,7,7,14,14,14,14,9,9,14,14,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,10,10,12,11,12,12,1,1,1,1,1,1,1,1,1,1,12,12,12,12,5,5,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,7,7,14,14,14,14,9,9,14,14,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,10,10,11,11,12,12,1,1,1,1,1,1,1,1,12,1,12,1,12,12,12,12,11,11,11,11,11,11,11,11,11,11,3,3,6,6,2,2,6,6,6,6,4,4,7,7,14,14,14,14,14,14,9,9,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,10,15,11,11,11,12,12,12,1,1,1,1,1,1,1,12,1,12,12,12,12,12,11,11,11,11,11,11,11,11,11,11,3,13,6,6,2,2,6,6,4,4,4,4,7,7,14,14,14,14,14,14,9,9,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,10,10,11,11,12,12,1,1,1,1,1,1,12,1,12,1,12,12,5,5,5,5,5,5,5,5,5,5,5,5,2,5,2,2,2,2,2,2,2,2,2,2,2,2,9,7,14,14,14,14,14,14,9,9,14,14,14,14,14,14,9,9,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,10,10,11,11,12,12,1,1,1,1,1,1,1,12,1,1,12,12,5,5,5,5,5,5,5,5,5,5,5,5,5,2,2,2,2,2,2,2,2,2,2,2,2,2,9,7,14,14,14,14,14,14,9,9,14,14,14,14,14,14,9,9,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,10,10,10,12,11,12,1,1,1,1,1,1,1,12,1,6,6,6,6,5,5,0,0,0,0,0,0,0,0,0,0,0,8,0,0,0,0,0,0,0,0,3,3,3,6,7,7,14,14,14,14,14,14,14,14,9,9,9,9,9,9,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,10,10,11,11,1,12,1,1,1,1,1,1,1,12,6,6,6,6,5,5,3,0,0,0,0,8,0,0,0,8,0,8,0,0,0,0,3,0,3,8,3,3,3,3,7,9,14,14,14,14,14,14,14,14,9,9,9,9,9,9,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,10,10,11,11,12,1,1,1,1,1,12,1,12,1,6,6,8,0,2,2,0,3,6,6,6,6,8,0,6,6,6,6,8,8,8,8,6,6,6,6,8,0,4,6,2,2,7,7,14,14,14,14,14,14,14,14,14,14,9,9,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,10,10,10,11,11,1,12,1,1,1,1,1,12,1,12,6,3,3,0,2,2,3,0,6,6,6,6,8,0,6,6,6,6,8,8,8,8,6,6,6,6,8,0,6,4,2,2,9,7,14,14,14,14,14,14,14,14,14,14,9,9,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,10,10,11,11,12,12,1,1,1,1,12,1,12,12,6,6,0,3,5,2,0,0,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,3,3,6,3,7,7,14,14,14,14,14,14,14,14,9,9,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,10,10,11,11,12,12,1,1,1,1,1,12,12,12,6,6,0,0,2,5,0,0,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,0,8,3,3,7,7,14,14,14,14,14,14,14,14,9,9,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,10,10,11,11,11,12,12,1,1,1,12,1,12,12,5,5,5,5,5,2,0,0,6,6,6,6,8,8,6,6,6,6,8,8,8,8,6,6,6,6,8,8,6,6,2,2,3,3,9,9,14,14,14,14,14,14,9,9,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,10,15,11,12,12,12,1,12,1,1,1,12,12,12,5,5,5,5,2,5,0,0,6,6,6,6,8,8,6,6,6,6,8,8,8,8,6,3,6,6,8,8,6,6,2,2,6,3,9,7,14,14,14,14,14,14,9,9,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,10,10,11,11,12,1,1,1,12,1,12,12,5,5,0,3,0,0,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,3,3,3,6,9,7,14,14,14,14,9,9,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,10,10,10,1,11,1,12,1,1,1,12,12,12,5,5,3,0,0,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,0,0,3,3,3,3,9,7,14,14,14,14,9,9,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,10,10,11,11,12,12,12,1,12,1,12,12,5,5,0,0,6,6,0,0,6,6,6,6,8,0,6,6,6,6,8,8,8,8,6,6,6,6,8,0,6,6,2,2,7,7,14,14,9,9,9,9,9,9,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,10,10,11,11,12,12,1,12,1,12,12,12,5,5,3,3,6,6,0,0,6,6,6,6,8,0,6,6,6,6,8,8,8,8,6,6,6,6,8,0,6,4,2,2,7,7,14,14,9,9,9,9,9,9,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,10,10,12,12,12,1,12,1,12,12,5,5,0,0,0,3,0,0,0,3,8,3,0,3,0,3,8,3,8,0,0,0,0,3,8,3,0,0,3,3,3,3,7,7,14,14,14,14,14,14,9,9,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,10,10,10,12,11,12,12,1,12,12,12,5,5,8,0,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,3,3,6,3,9,7,14,14,14,14,14,14,9,9,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,10,2,11,12,12,1,12,1,12,12,5,5,5,5,5,5,5,5,2,2,2,2,2,2,2,2,2,2,5,2,5,2,5,2,2,2,2,2,2,2,7,7,14,14,14,14,14,14,9,9,9,9,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,10,10,12,11,12,12,1,12,12,12,5,5,5,5,5,5,5,5,2,2,2,2,2,2,2,2,2,2,2,5,2,5,2,5,2,2,2,2,2,2,7,7,14,14,14,14,14,14,9,9,9,9,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,10,10,10,10,1,12,1,1,1,1,12,1,12,1,12,12,12,12,11,12,2,2,6,6,2,2,6,6,6,6,6,6,6,6,6,6,6,6,6,4,4,4,7,7,14,14,14,14,14,14,9,9,14,14,9,9,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,10,10,10,10,2,12,12,12,12,1,1,1,12,12,12,12,12,12,12,12,11,2,2,6,6,2,2,6,6,6,6,6,6,6,6,6,6,6,6,4,6,4,4,7,7,14,14,14,14,14,14,9,9,14,14,9,9,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,10,10,11,11,12,11,12,1,1,1,1,1,1,1,12,1,12,1,12,12,12,12,5,5,3,3,2,2,3,0,3,3,0,0,0,0,0,0,0,0,3,3,3,6,7,7,14,14,14,14,9,9,14,14,14,14,9,9,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,10,10,10,11,11,11,12,12,12,12,12,1,1,1,1,1,12,1,12,12,12,12,12,5,2,0,3,2,2,0,3,0,0,8,8,0,8,0,0,0,8,3,0,3,3,7,7,14,14,14,14,9,9,14,14,14,14,9,9,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,10,10,12,11,12,12,12,12,12,1,1,1,1,1,1,1,1,1,1,1,12,1,12,12,5,5,5,2,2,5,3,0,0,0,6,6,6,6,8,8,6,6,6,6,3,3,7,7,14,14,14,14,9,9,14,14,14,14,14,14,9,9,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,10,10,10,11,11,11,12,12,1,1,12,1,1,1,1,1,1,1,1,1,1,1,12,12,12,5,5,5,5,5,2,0,0,0,0,6,6,6,6,8,8,6,6,6,6,3,3,7,7,14,14,14,14,9,9,14,14,14,14,14,14,9,9,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,10,10,12,11,12,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,1,12,12,11,12,5,5,0,0,8,8,8,8,8,8,8,8,8,8,8,8,3,3,3,6,7,7,14,14,9,9,14,14,14,14,14,14,9,9,9,9,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,10,10,11,11,12,12,1,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,12,12,12,11,5,5,0,0,8,8,8,8,8,8,8,8,8,8,8,8,3,3,3,3,7,7,14,14,9,9,14,14,14,14,14,14,9,9,9,9,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,15,10,10,11,11,12,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,1,12,12,5,5,0,0,0,0,6,6,6,6,8,0,6,6,6,6,8,3,4,6,7,7,14,14,9,9,14,14,9,9,9,9,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,15,10,10,11,11,11,12,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,12,12,5,5,0,0,0,0,6,6,6,6,8,0,6,6,6,6,3,8,4,4,7,7,14,14,9,9,14,14,9,9,9,9,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,10,10,10,12,11,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,1,12,12,5,5,0,0,0,3,8,0,8,0,8,0,8,0,8,0,0,3,3,3,3,3,7,9,14,14,9,9,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,15,10,10,12,11,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,12,12,5,5,8,0,3,0,8,0,0,0,0,0,0,0,0,0,3,0,3,3,3,6,9,7,14,14,9,9,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,10,10,11,11,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,1,12,12,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,2,2,2,7,7,14,14,9,9,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,10,10,10,11,11,12,12,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,12,12,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,2,2,2,2,7,9,14,14,9,9,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,10,10,12,11,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,1,12,1,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,0,3,3,2,2,9,7,14,14,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,10,10,12,11,1,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,0,13,3,0,2,2,9,7,14,14,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,10,10,11,11,12,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,1,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,0,8,6,3,9,7,14,14,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,10,15,11,11,11,12,1,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,3,0,3,8,7,7,14,14,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,10,10,11,11,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,1,12,1,12,1,12,1,12,1,12,13,13,13,13,13,13,8,8,7,7,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,10,10,11,11,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,1,12,1,12,1,12,1,12,1,12,1,12,1,13,13,13,13,13,13,0,0,7,7,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,10,10,10,12,11,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,3,0,7,7,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,10,10,11,11,1,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,0,3,7,7,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,10,10,11,11,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,8,0,3,3,7,7,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,10,10,10,11,11,1,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,3,0,7,7,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,10,10,11,11,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,0,3,7,7,7,7,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,10,10,11,11,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,1,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,3,0,7,7,7,7,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,10,10,11,11,11,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,13,13,13,13,13,13,13,13,13,13,13,13,13,13,8,13,13,0,13,13,8,0,3,8,3,3,7,7,14,14,9,9,14,14,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,10,15,11,12,12,12,1,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,1,13,13,13,13,13,13,13,13,13,13,13,13,0,13,13,8,13,13,0,13,13,13,13,3,3,0,7,7,14,14,9,9,14,14,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,10,10,12,11,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,13,13,13,13,13,13,13,13,13,13,5,5,5,5,5,5,2,5,2,5,5,5,2,2,2,2,7,7,14,14,14,14,9,9,14,14,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,10,10,10,12,11,1,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,13,13,13,13,13,13,13,13,13,13,2,5,5,5,5,5,5,5,5,5,5,5,2,2,2,2,7,7,14,14,14,14,9,9,14,14,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,10,10,11,11,11,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,13,13,13,13,13,13,13,13,8,13,5,5,0,0,6,6,6,6,0,3,6,6,6,6,3,3,7,7,14,14,14,14,14,14,9,9,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,10,10,11,12,12,12,1,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,13,13,13,13,13,13,13,13,13,3,5,5,3,3,6,6,6,6,3,0,6,6,6,4,3,6,7,7,14,14,14,14,14,14,9,9,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,15,10,10,12,11,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,13,13,13,13,13,13,8,0,13,13,5,5,0,0,0,0,0,0,8,0,0,0,3,3,3,3,7,7,14,14,14,14,14,14,9,9,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,10,10,10,12,11,1,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,13,13,13,13,13,13,13,13,0,13,2,2,3,0,0,8,0,8,0,0,0,8,3,0,3,3,7,7,14,14,14,14,14,14,9,9,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,15,10,10,11,11,12,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,13,13,13,13,5,5,2,5,2,2,5,5,0,3,6,6,6,6,8,8,6,6,6,6,3,3,7,7,14,14,14,14,14,14,14,14,9,9,9,9,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,15,10,10,11,11,11,12,1,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,13,13,13,13,5,5,5,5,5,5,2,2,3,0,6,6,6,6,8,8,6,6,6,6,3,3,7,7,14,14,14,14,14,14,14,14,9,9,9,9,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,10,10,11,11,12,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,13,13,13,13,5,5,0,0,3,3,2,5,0,0,8,0,8,8,8,8,8,0,8,0,3,3,3,6,7,7,14,14,14,14,14,14,14,14,14,14,9,9,9,9,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,10,10,11,12,12,12,1,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,13,13,13,13,5,5,3,3,0,0,2,2,0,0,0,8,8,8,8,8,8,0,0,0,3,3,3,3,9,7,14,14,14,14,14,14,14,14,14,14,9,9,9,9,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,10,15,10,10,11,11,12,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,12,5,5,0,0,6,6,5,5,0,0,6,6,6,6,0,3,6,6,6,6,3,3,4,4,7,7,14,14,14,14,14,14,14,14,14,14,9,9,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,10,10,1,12,12,12,1,12,1,1,1,1,1,1,1,1,1,1,1,1,12,12,12,12,5,5,3,0,6,6,2,2,3,3,6,6,6,6,0,0,6,6,6,6,3,3,4,4,9,7,14,14,14,14,14,14,14,14,14,14,9,9,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,10,15,10,10,1,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,12,5,5,0,3,0,0,5,5,0,0,0,0,8,0,5,2,5,2,2,2,2,2,2,2,9,7,9,9,14,14,14,14,14,14,9,9,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,10,10,2,12,12,1,12,1,1,1,1,1,1,1,1,1,1,1,1,12,12,12,12,5,5,3,0,3,0,2,2,3,3,0,3,0,3,2,5,2,5,2,2,2,2,2,2,9,9,9,9,14,14,14,14,14,14,9,9,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,10,10,10,10,12,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,12,5,5,0,0,3,3,2,2,6,6,6,6,6,6,2,2,3,3,3,0,3,3,4,3,9,7,9,9,14,14,14,14,14,14,9,9,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,10,10,10,1,12,1,12,1,1,1,1,1,1,1,1,1,1,1,1,12,12,12,12,5,5,3,3,0,3,2,2,6,4,6,6,6,6,2,2,0,0,3,3,3,3,3,3,9,7,9,9,14,14,14,14,14,14,9,9,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,10,10,1,11,1,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,12,5,5,6,6,6,6,2,2,6,6,6,6,4,6,2,2,3,3,6,6,4,6,7,7,14,14,14,14,9,9,9,9,9,9,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,10,10,12,11,12,12,1,12,1,1,1,1,1,1,1,1,1,1,1,1,12,12,12,12,5,5,6,6,6,6,2,2,6,6,4,6,6,6,2,2,3,0,6,6,4,4,7,7,14,14,14,14,9,9,9,9,9,9,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,10,10,11,11,12,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,12,5,5,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,6,7,7,14,14,14,14,14,14,14,14,9,9,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,10,10,11,11,11,12,1,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,12,12,12,5,5,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,7,7,14,14,14,14,14,14,14,14,9,9,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,15,15,10,10,10,12,11,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,1,12,1,12,12,12,12,11,11,11,11,11,11,11,11,11,11,3,3,6,6,2,2,6,6,6,4,4,4,7,7,14,14,14,14,14,14,14,14,9,9,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,10,10,12,11,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,12,1,12,12,12,12,12,11,11,11,11,11,11,11,11,11,11,3,13,6,6,2,2,6,6,4,6,4,4,7,7,14,14,14,14,14,14,14,14,9,9,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,15,10,10,11,11,12,12,1,1,1,1,1,1,1,1,1,1,1,1,12,1,12,1,12,12,5,5,5,5,5,5,5,5,5,5,5,5,2,5,2,2,2,2,2,2,2,2,2,2,2,2,7,7,14,14,14,14,14,14,9,9,9,9,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,10,10,10,11,11,12,12,12,12,1,1,1,1,1,1,1,1,1,1,1,12,1,1,12,12,5,5,5,5,5,5,5,5,5,5,5,5,5,2,2,2,2,2,2,2,2,2,2,2,2,2,7,7,14,14,14,14,14,14,9,9,9,9,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,15,10,10,12,11,12,1,1,1,1,1,1,1,1,1,1,1,1,1,12,1,6,6,6,6,5,5,0,0,0,0,0,0,0,0,0,0,0,8,0,0,0,0,0,0,0,0,3,3,3,3,3,6,7,7,14,14,14,14,9,9,14,14,9,9,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,15,10,10,12,11,1,12,1,1,1,1,1,1,1,1,1,1,1,1,1,12,6,6,6,6,5,5,3,0,0,0,0,8,0,0,0,8,0,8,0,0,0,0,3,0,3,8,0,0,3,3,3,3,7,7,14,14,14,14,9,9,14,14,9,9,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,10,10,11,11,12,12,12,1,1,1,1,1,1,1,1,1,1,1,12,1,12,1,6,6,8,0,2,2,0,3,6,6,6,6,8,0,6,6,6,6,8,8,8,8,6,6,6,6,0,0,6,6,4,4,7,7,14,14,9,9,14,14,14,14,9,9,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,10,15,11,11,11,12,1,12,1,1,1,1,1,1,1,1,1,1,1,12,1,12,6,3,3,0,2,2,3,0,6,6,6,6,8,0,6,6,6,6,8,8,8,8,6,6,6,6,8,0,6,6,4,6,7,7,14,14,7,9,14,14,14,14,9,9,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,10,10,11,11,12,12,1,1,1,1,1,1,1,1,1,1,1,1,12,1,12,12,6,6,0,3,5,2,0,0,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,0,3,3,3,7,9,9,9,14,14,14,14,14,14,9,9,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,10,10,11,11,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,12,12,12,6,6,0,0,2,5,0,0,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,3,0,3,6,7,7,9,9,14,14,14,14,14,14,9,9,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,10,10,10,12,11,12,1,1,1,1,1,1,1,1,1,1,1,1,1,12,1,12,12,5,5,5,5,5,2,0,0,6,6,6,6,8,8,6,6,6,6,8,8,8,8,6,6,6,6,8,8,6,6,6,6,3,3,7,7,7,7,14,14,14,14,14,14,9,9,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,10,10,11,11,1,12,1,1,1,1,1,1,1,1,1,1,1,1,1,12,12,12,5,5,5,5,2,5,0,0,6,6,6,6,8,8,6,6,6,6,8,8,8,8,6,3,6,6,8,8,6,6,6,6,3,3,7,7,9,9,14,14,14,14,14,14,9,9,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,10,10,11,11,12,1,1,1,1,1,1,1,1,1,1,1,1,1,12,1,12,12,5,5,0,3,0,0,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,0,3,3,3,3,9,7,14,14,14,14,14,14,14,14,9,9,14,14,14),
(15,15,15,15,15,15,15,15,15,15,10,10,10,11,11,1,12,1,1,1,1,1,1,1,1,1,1,1,1,1,12,12,12,5,5,3,0,0,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,3,3,3,4,7,9,14,14,14,14,14,14,14,14,9,9,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,10,10,11,11,12,12,1,1,1,1,1,1,1,1,1,1,1,1,12,1,12,12,5,5,0,0,6,6,0,0,6,6,6,6,8,0,6,6,6,6,8,8,8,8,6,6,6,6,8,0,6,6,6,6,3,3,2,2,9,7,14,14,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,10,10,11,11,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,12,12,12,5,5,3,3,6,6,0,0,6,6,6,6,8,0,6,6,6,6,8,8,8,8,6,6,6,6,8,0,6,6,6,6,3,3,2,2,9,7,14,14,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,10,10,11,11,11,12,12,1,1,1,1,1,1,1,1,1,1,1,12,1,12,12,5,5,0,0,0,3,0,0,0,3,8,3,0,3,0,3,8,3,8,0,0,0,0,3,8,3,0,3,0,3,3,3,3,6,7,7,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,10,10,11,11,12,12,1,12,1,1,1,1,1,1,1,1,1,1,1,12,12,12,5,5,8,0,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,3,3,7,7,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,15,10,10,12,11,12,1,1,1,1,1,1,1,1,1,1,1,12,1,12,12,5,5,5,5,5,5,5,5,2,2,2,2,2,2,2,2,2,2,5,2,5,2,5,2,2,2,2,2,2,2,2,2,2,2,7,7,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,15,10,2,12,11,1,12,1,1,1,1,1,1,1,1,1,1,1,12,12,12,5,5,5,5,5,5,5,5,2,2,2,2,2,2,2,2,2,2,2,5,2,5,2,5,2,2,2,2,2,2,2,2,2,2,7,7,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,10,10,10,10,12,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,12,1,12,1,12,12,12,12,11,12,2,2,6,6,2,2,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,4,4,4,4,7,7,14,14,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,10,10,10,1,12,1,12,1,1,1,1,1,1,1,1,1,1,1,1,1,12,12,12,12,12,12,12,12,11,2,2,6,6,2,2,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,4,6,4,4,9,7,14,14,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,10,10,1,11,1,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,1,12,1,12,12,12,12,5,5,3,3,2,2,3,0,3,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,3,3,7,7,14,14,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,10,10,12,11,12,12,1,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,1,12,12,12,12,12,5,2,0,3,2,2,0,3,0,0,8,8,0,8,0,0,0,8,0,8,0,0,0,8,3,0,3,6,7,7,14,14,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,10,10,11,11,12,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,1,12,12,5,5,5,2,2,5,3,0,0,0,6,6,6,6,8,8,6,6,6,6,8,8,6,6,6,6,3,3,7,7,14,14,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,10,10,11,11,11,12,1,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,12,12,5,5,5,5,5,2,0,0,0,0,6,6,6,6,8,8,6,6,6,6,8,8,6,6,6,6,3,3,7,7,14,14,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,10,10,10,12,11,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,1,12,12,11,12,5,5,0,0,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,0,3,3,3,3,9,7,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,10,10,12,11,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,12,12,12,11,5,5,0,0,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,3,3,6,3,9,9,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,10,10,11,11,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,1,12,12,5,5,0,0,0,0,6,6,6,6,8,0,6,6,6,6,8,0,6,6,6,4,3,3,7,7,9,9,14,14,14,14,14,14,9,9,14,14,14),
(15,15,15,15,15,15,10,10,10,11,11,12,12,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,12,12,5,5,0,0,0,0,6,6,6,6,8,0,6,6,6,6,8,0,6,6,6,4,3,3,7,7,9,7,14,14,14,14,14,14,9,9,14,14,14),
(15,15,15,15,15,15,15,10,10,12,11,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,1,12,12,5,5,0,0,0,3,8,0,8,0,8,0,8,0,8,0,8,0,3,3,3,0,7,7,14,14,14,14,9,9,14,14,9,9,14,14,14,14,14),
(15,15,15,15,15,15,15,10,10,12,11,1,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,12,12,5,5,8,0,3,0,8,0,0,0,0,0,0,0,0,0,0,0,3,3,3,4,7,7,14,14,14,14,9,9,14,14,9,9,14,14,14,14,14),
(15,15,15,15,15,10,10,11,11,12,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,1,12,12,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,2,2,2,2,9,7,14,14,14,14,9,9,14,14,9,9,14,14,14,14,14),
(15,15,15,15,15,10,15,11,11,11,12,1,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,12,12,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,2,5,2,2,2,2,7,7,14,14,14,14,9,9,14,14,9,9,14,14,14,14,14),
(15,15,15,15,15,10,10,11,11,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,1,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,8,13,0,3,0,7,7,14,14,14,14,14,14,14,14,9,9,14,14,14,14,14,14,14),
(15,15,15,15,15,10,10,11,11,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,3,3,7,7,14,14,14,14,14,14,14,14,9,9,14,14,14,14,14,14,14),
(15,15,15,15,10,10,10,12,11,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,1,13,13,13,13,13,13,13,13,13,13,13,13,13,13,0,0,3,3,7,7,14,14,14,14,14,14,14,14,9,9,14,14,14,14,14,14,14),
(15,15,15,15,15,10,10,11,11,1,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,3,0,7,7,14,14,14,14,14,14,14,14,9,9,14,14,14,14,14,14,14),
(15,15,15,15,15,10,10,11,11,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,13,13,13,13,13,13,13,13,13,13,13,13,13,13,0,0,7,7,14,14,14,14,14,14,14,14,9,9,14,14,14,14,14,14,14,14,14),
(15,15,15,15,10,10,10,11,11,1,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,1,13,13,13,13,13,13,13,13,13,13,13,13,13,13,8,0,7,7,14,14,14,14,14,14,14,14,9,9,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,10,10,11,11,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,1,12,1,12,1,12,1,12,1,12,13,13,0,0,7,7,14,14,14,14,14,14,14,14,9,9,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,10,10,11,11,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,1,12,1,1,1,1,1,1,1,1,1,1,1,13,13,0,3,7,7,14,14,14,14,14,14,14,14,9,9,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,10,10,11,11,11,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,0,0,7,7,14,14,14,14,14,14,14,14,9,9,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,10,15,11,12,12,12,1,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,0,3,7,7,14,14,14,14,14,14,14,14,9,9,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,10,10,12,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,8,8,7,7,14,14,14,14,14,14,14,14,9,9,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,10,10,10,1,11,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,8,3,7,7,14,14,14,14,14,14,14,14,9,9,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,10,10,12,11,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,8,13,3,0,7,7,14,14,14,14,14,14,14,14,9,9,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,10,10,12,11,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,1,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,3,3,3,7,7,14,14,14,14,14,14,14,14,9,9,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,10,15,11,11,12,12,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,13,13,13,13,13,13,13,13,13,13,13,13,13,13,8,13,13,0,13,13,0,0,13,3,3,3,7,7,14,14,14,14,14,14,9,9,9,9,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,10,10,11,12,11,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,1,13,13,13,13,13,13,13,13,13,13,13,13,0,13,13,8,13,13,0,13,13,13,0,13,3,3,7,7,14,14,14,14,14,14,9,9,9,9,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,10,10,12,11,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,13,13,13,13,13,13,13,13,13,13,5,5,5,5,5,5,2,5,2,5,5,5,2,5,5,2,2,2,2,2,9,7,14,14,9,9,14,14,14,14,9,9,14,14,14,14,14),
(15,15,15,15,15,15,15,15,10,10,10,12,11,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,13,13,13,13,13,13,13,13,13,13,2,5,5,5,5,5,5,5,5,5,5,5,5,5,2,2,2,2,2,2,9,7,14,14,9,9,14,14,14,14,9,9,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,10,10,11,11,11,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,13,13,13,13,13,13,13,13,8,13,5,5,0,0,6,6,6,6,0,3,6,6,6,6,0,3,6,4,4,4,7,7,14,14,9,9,14,14,14,14,9,9,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,10,10,11,12,12,12,1,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,13,13,13,13,13,13,13,13,13,3,5,5,3,3,6,6,6,6,3,0,6,6,6,6,3,0,4,6,4,4,7,7,14,14,9,9,14,14,14,14,9,9,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,10,10,12,11,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,13,13,13,13,13,13,8,0,13,13,5,5,0,0,0,0,0,0,8,0,0,0,8,0,8,0,0,0,3,3,3,6,7,9,14,14,14,14,14,14,14,14,9,9,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,10,10,12,11,1,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,13,13,13,13,13,13,13,13,0,13,2,2,3,0,0,8,0,8,0,0,0,8,0,8,0,0,0,8,3,3,3,3,9,7,14,14,14,14,14,14,14,14,9,9,14,14,14),
(15,15,15,15,15,15,15,15,15,15,10,10,10,12,11,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,13,13,13,13,5,5,2,5,2,2,5,5,0,3,6,6,6,6,8,8,6,6,6,6,8,8,6,6,6,6,3,6,7,7,14,14,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,10,10,12,12,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,13,13,13,13,5,5,5,5,5,5,2,2,3,0,6,6,6,6,8,8,6,6,6,6,8,8,6,6,4,4,3,3,9,7,14,14,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,10,10,10,10,1,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,13,13,13,13,5,5,0,0,3,3,2,5,0,0,8,0,8,8,8,8,8,0,8,0,8,0,8,3,0,3,7,7,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,10,10,10,10,2,12,12,1,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,13,13,13,13,5,5,3,3,0,0,2,2,0,0,0,8,8,8,8,8,8,0,0,0,0,0,3,3,3,3,7,7,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,10,10,1,11,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,12,5,5,0,0,6,6,5,5,0,0,6,6,6,6,0,3,6,6,6,6,0,3,6,6,4,4,9,7,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,10,10,10,12,11,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,12,12,12,5,5,3,0,6,6,2,2,3,3,6,6,6,6,0,0,6,6,6,6,3,0,4,4,4,4,7,7,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,10,10,12,11,12,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,12,5,5,0,3,0,0,5,5,0,0,0,0,8,0,5,2,5,2,5,2,2,2,2,2,2,2,9,9,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,10,10,10,12,11,12,12,1,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,12,12,12,5,5,3,0,3,0,2,2,3,3,0,3,0,3,2,5,2,5,2,5,2,2,2,2,2,2,9,7,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,10,10,12,11,12,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,12,5,5,0,0,3,3,2,2,6,6,6,6,6,6,2,2,3,3,0,3,3,3,3,6,9,7,9,9,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,10,10,11,11,11,12,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,12,12,12,5,5,3,3,0,3,2,2,6,4,6,6,6,6,2,2,0,0,3,0,3,0,3,3,7,7,9,7,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,10,10,11,11,12,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,12,5,5,6,6,6,6,2,2,6,6,6,6,4,6,2,2,3,3,6,6,4,4,3,6,7,7,14,14,9,9,14,14,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,10,10,11,11,11,12,1,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,12,12,12,5,5,6,6,6,6,2,2,6,6,4,6,6,6,2,2,3,0,6,6,6,4,3,3,9,7,14,14,9,9,14,14,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,10,10,10,12,11,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,12,5,5,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,7,7,14,14,14,14,9,9,14,14,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,10,10,12,11,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,12,12,12,5,5,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,6,7,7,14,14,14,14,9,9,14,14,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,10,10,11,11,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,1,12,1,12,12,12,12,11,11,11,11,11,11,11,11,11,11,3,3,6,6,2,2,6,6,6,6,4,4,7,7,14,14,14,14,14,14,9,9,14,14,14,14,14,14,14,14,14,14,14),
(15,15,10,10,10,11,11,12,12,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,1,12,12,12,12,12,11,11,11,11,11,11,11,11,11,11,3,13,6,6,2,2,6,6,4,6,4,4,7,7,14,14,14,14,14,14,9,9,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,10,10,12,11,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,1,12,1,12,12,5,5,5,5,5,5,5,5,5,5,5,5,2,5,2,2,2,2,2,2,2,2,2,2,2,2,9,7,14,14,14,14,14,14,9,9,14,14,14,14,14,14,9,9,14,14,14),
(15,15,15,10,10,12,11,1,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,1,1,12,12,5,5,5,5,5,5,5,5,5,5,5,5,5,2,2,2,2,2,2,2,2,2,2,2,2,2,9,7,14,14,14,14,14,14,9,9,14,14,14,14,14,14,9,9,14,14,14),
(15,10,10,11,11,12,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,1,6,6,6,6,5,5,0,0,0,0,0,0,0,0,0,0,0,8,0,0,0,0,0,0,0,0,3,3,3,6,7,7,14,14,14,14,14,14,14,14,9,9,9,9,9,9,14,14,14,14,14),
(15,10,15,11,11,11,12,1,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,6,6,6,6,5,5,3,0,0,0,0,8,0,0,0,8,0,8,0,0,0,0,3,0,3,8,3,3,3,3,7,7,14,14,14,14,14,14,14,14,9,9,9,9,9,9,14,14,14,14,14),
(15,10,10,11,11,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,1,12,1,6,6,8,0,2,2,0,3,6,6,6,6,8,0,6,6,6,6,8,8,8,8,6,6,6,6,8,0,4,4,4,4,7,9,14,14,14,14,14,14,14,14,14,14,9,9,14,14,14,14,14),
(15,10,10,11,11,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,1,12,6,3,3,0,2,2,3,0,6,6,6,6,8,0,6,6,6,6,8,8,8,8,6,6,6,6,8,0,4,6,4,4,7,7,14,14,14,14,14,14,14,14,14,14,9,9,14,14,14,14,14),
(15,10,10,12,11,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,1,12,12,6,6,0,3,5,2,0,0,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,0,3,3,7,7,14,14,14,14,14,14,14,14,9,9,14,14,14,14,14,14,14),
(15,10,10,12,11,1,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,12,12,6,6,0,0,2,5,0,0,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,0,8,3,3,7,7,14,14,14,14,14,14,14,14,9,9,14,14,14,14,14,14,14),
(15,10,10,11,11,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,1,12,12,5,5,5,5,5,2,0,0,6,6,6,6,8,8,6,6,6,6,8,8,8,8,6,6,6,6,8,8,6,6,4,6,3,3,7,9,14,14,14,14,14,14,9,9,14,14,14,14,14,14,14),
(15,10,10,12,11,1,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,12,12,5,5,5,5,2,5,0,0,6,6,6,6,8,8,6,6,6,6,8,8,8,8,6,3,6,6,8,8,6,6,6,4,3,3,9,7,14,14,14,14,14,14,9,9,14,14,14,14,14,14,14),
(15,10,10,11,11,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,1,12,12,5,5,0,3,0,0,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,0,3,0,3,6,9,7,14,14,14,14,9,9,14,14,14,14,14,14,14,14,14),
(15,10,10,11,11,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,12,12,5,5,3,0,0,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,0,0,3,3,3,3,7,7,14,14,14,14,9,9,14,14,14,14,14,14,14,14,14),
(15,10,10,11,11,11,12,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,1,12,12,5,5,0,0,6,6,0,0,6,6,6,6,8,0,6,6,6,6,8,8,8,8,6,6,6,6,8,0,6,6,4,4,7,7,14,14,9,9,9,9,9,9,14,14,14,14,14,14,14,14,14),
(15,10,15,11,12,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,12,12,5,5,3,3,6,6,0,0,6,6,6,6,8,0,6,6,6,6,8,8,8,8,6,6,6,6,8,0,6,6,4,4,7,7,14,14,7,9,9,9,9,9,14,14,14,14,14,14,14,14,14),
(15,15,15,10,10,12,11,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,1,12,12,5,5,0,0,0,3,0,0,0,3,8,3,0,3,0,3,8,3,8,0,0,0,0,3,8,3,0,3,3,3,3,6,7,7,14,14,14,14,14,14,9,9,14,14,14,14,14,14,14,14,14),
(15,15,10,10,10,12,11,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,12,12,5,5,8,0,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,3,3,7,7,14,14,14,14,14,14,9,9,14,14,14,14,14,14,14,14,14),
(15,15,15,10,10,11,11,11,12,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,1,12,12,5,5,5,5,5,5,5,5,2,2,2,2,2,2,2,2,2,2,5,2,5,2,5,2,2,2,2,2,2,2,7,7,14,14,14,14,14,14,9,9,9,9,14,14,14,14,14,14,14,14,14),
(15,15,15,10,10,11,12,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,12,12,5,5,5,5,5,5,5,5,2,2,2,2,2,2,2,2,2,2,2,5,2,5,2,5,2,2,2,2,2,2,7,7,14,14,14,14,14,14,9,9,9,9,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,10,10,11,11,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,1,12,1,12,12,12,12,11,12,2,2,6,6,2,2,6,6,6,6,6,6,6,6,6,6,6,6,6,4,4,4,7,7,14,14,14,14,14,14,9,9,14,14,9,9,14,14,14,14,14,14,14),
(15,15,15,15,10,10,10,12,11,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,12,12,12,12,12,12,12,11,2,2,6,6,2,2,6,6,6,6,6,6,6,6,6,6,6,6,4,6,4,4,7,7,14,14,14,14,14,14,9,9,14,14,9,9,14,14,14,14,14,14,14),
(15,15,15,15,15,10,10,11,11,11,11,1,1,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,1,12,1,12,12,12,12,5,5,3,3,2,2,3,0,3,3,0,0,0,0,0,0,0,0,3,3,3,6,7,7,14,14,14,14,9,9,14,14,14,14,9,9,14,14,14,14,14,14,14),
(15,15,15,15,15,10,10,11,11,12,11,12,12,1,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,1,12,12,12,12,12,5,2,0,3,2,2,0,3,0,0,8,8,0,8,0,0,0,8,3,0,3,3,7,7,14,14,14,14,9,9,14,14,14,14,9,9,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,10,10,11,11,11,11,12,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,1,12,12,5,5,5,2,2,5,3,0,0,0,6,6,6,6,8,8,6,6,6,6,3,3,7,7,14,14,14,14,9,9,14,14,14,14,14,14,9,9,14,14,14,14,14),
(15,15,15,15,15,15,15,10,10,11,11,11,1,12,12,1,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,12,12,5,5,5,5,5,2,0,0,0,0,6,6,6,6,8,8,6,6,6,6,3,3,7,7,14,14,14,14,9,9,14,14,14,14,14,14,9,9,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,10,10,10,10,12,11,12,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,1,12,12,11,12,5,5,0,0,8,8,8,8,8,8,8,8,8,8,8,8,3,3,3,6,7,7,14,14,9,9,14,14,14,14,14,14,9,9,9,9,14,14,14),
(15,15,15,15,15,15,15,15,15,10,10,10,10,1,11,12,12,1,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,12,12,12,11,5,5,0,0,8,8,8,8,8,8,8,8,8,8,8,8,3,3,3,3,7,7,14,14,9,9,14,14,14,14,14,14,9,9,9,9,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,10,10,10,2,11,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,1,12,12,5,5,0,0,0,0,6,6,6,6,8,0,6,6,6,6,8,3,4,6,7,7,14,14,9,9,14,14,9,9,9,9,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,10,10,10,10,1,12,1,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,12,12,5,5,0,0,0,0,6,6,6,6,8,0,6,6,6,6,3,8,4,4,7,7,14,14,9,9,14,14,9,9,9,9,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,10,10,10,1,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,1,12,12,5,5,0,0,0,3,8,0,8,0,8,0,8,0,8,0,0,3,3,3,3,3,7,9,14,14,9,9,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,15,10,10,1,11,1,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,12,12,5,5,8,0,3,0,8,0,0,0,0,0,0,0,0,0,3,0,3,3,3,6,9,7,14,14,9,9,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,10,10,11,11,12,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,1,12,12,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,2,2,2,7,7,14,14,9,9,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,10,10,10,11,11,12,12,1,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,12,12,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,2,2,2,2,7,9,14,14,9,9,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,10,10,12,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,1,12,1,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,0,3,3,2,2,9,7,14,14,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,10,10,12,11,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,0,13,3,0,2,2,9,7,14,14,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,10,10,11,11,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,1,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,0,8,6,3,9,7,14,14,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,10,15,11,11,11,12,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,3,0,3,8,7,7,14,14,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,10,10,11,11,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,1,12,1,12,1,12,1,12,1,12,13,13,13,13,13,13,8,8,7,7,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,10,10,11,11,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,1,12,1,12,1,12,1,12,1,12,1,12,1,13,13,13,13,13,13,0,0,7,7,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,10,10,10,12,11,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,3,0,7,7,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,10,10,11,11,1,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,0,3,7,7,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,10,10,11,11,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,8,0,3,3,7,7,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,10,10,10,11,11,1,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,3,0,7,7,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,10,10,11,11,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,0,3,7,7,7,7,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,10,10,11,11,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,1,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,3,0,7,7,7,7,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,10,10,11,11,11,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,13,13,13,13,13,13,13,13,13,13,13,13,13,13,8,13,13,0,13,13,8,0,3,8,3,3,7,7,14,14,9,9,14,14,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,10,15,11,12,12,12,1,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,1,13,13,13,13,13,13,13,13,13,13,13,13,0,13,13,8,13,13,0,13,13,13,13,3,3,0,7,7,14,14,9,9,14,14,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,10,10,12,11,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,13,13,13,13,13,13,13,13,13,13,5,5,5,5,5,5,2,5,2,5,5,5,2,2,2,2,7,7,14,14,14,14,9,9,14,14,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,10,10,10,12,11,1,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,13,13,13,13,13,13,13,13,13,13,2,5,5,5,5,5,5,5,5,5,5,5,2,2,2,2,7,7,14,14,14,14,9,9,14,14,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,10,10,11,11,11,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,13,13,13,13,13,13,13,13,8,13,5,5,0,0,6,6,6,6,0,3,6,6,6,6,3,3,7,7,14,14,14,14,14,14,9,9,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,10,10,11,12,12,12,1,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,13,13,13,13,13,13,13,13,13,3,5,5,3,3,6,6,6,6,3,0,6,6,6,4,3,6,7,7,14,14,14,14,14,14,9,9,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,15,10,10,12,11,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,13,13,13,13,13,13,8,0,13,13,5,5,0,0,0,0,0,0,8,0,0,0,3,3,3,3,7,7,14,14,14,14,14,14,9,9,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,10,10,10,12,11,1,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,13,13,13,13,13,13,13,13,0,13,2,2,3,0,0,8,0,8,0,0,0,8,3,0,3,3,7,7,14,14,14,14,14,14,9,9,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,15,10,10,11,11,12,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,13,13,13,13,5,5,2,5,2,2,5,5,0,3,6,6,6,6,8,8,6,6,6,6,3,3,7,7,14,14,14,14,14,14,14,14,9,9,9,9,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,15,10,10,11,11,11,12,1,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,13,13,13,13,5,5,5,5,5,5,2,2,3,0,6,6,6,6,8,8,6,6,6,6,3,3,7,7,14,14,14,14,14,14,14,14,9,9,9,9,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,10,10,11,11,12,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,13,13,13,13,5,5,0,0,3,3,2,5,0,0,8,0,8,8,8,8,8,0,8,0,3,3,3,3,7,9,14,14,14,14,14,14,14,14,14,14,9,9,9,9,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,10,10,11,12,12,12,1,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,13,13,13,13,5,5,3,3,0,0,2,2,0,0,0,8,8,8,8,8,8,0,0,0,3,3,3,4,9,7,14,14,14,14,14,14,14,14,14,14,9,9,9,9,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,10,15,10,10,11,11,12,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,12,5,5,0,0,6,6,5,5,0,0,6,6,6,6,0,3,6,6,6,6,3,3,2,2,9,7,14,14,14,14,14,14,14,14,14,14,9,9,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,10,10,1,12,12,12,1,12,1,1,1,1,1,1,1,1,1,1,1,1,12,12,12,12,5,5,3,0,6,6,2,2,3,3,6,6,6,6,0,0,6,6,6,6,3,3,2,2,9,7,14,14,14,14,14,14,14,14,14,14,9,9,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,10,15,10,10,1,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,12,5,5,0,3,0,0,5,5,0,0,0,0,8,0,5,2,5,2,2,2,2,2,2,10,7,9,9,9,14,14,14,14,14,14,9,9,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,10,10,2,12,12,1,12,1,1,1,1,1,1,1,1,1,1,1,1,12,12,12,12,5,5,3,0,3,0,2,2,3,3,0,3,0,3,2,5,2,5,2,2,2,2,2,2,9,7,9,7,14,14,14,14,14,14,9,9,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,10,10,10,10,12,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,12,5,5,0,0,3,3,2,2,6,6,6,6,6,6,2,2,3,3,3,3,3,3,4,3,9,7,9,9,14,14,14,14,14,14,9,9,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,10,10,10,1,12,1,12,1,1,1,1,1,1,1,1,1,1,1,1,12,12,12,12,5,5,3,3,0,3,2,2,6,4,6,6,6,6,2,2,0,0,3,0,3,3,3,3,7,7,9,9,14,14,14,14,14,14,9,9,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,10,10,1,11,1,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,12,5,5,6,6,6,6,2,2,6,6,6,6,4,6,2,2,3,3,6,6,4,4,7,7,14,14,14,14,9,9,9,9,9,9,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,10,10,12,11,12,12,1,12,1,1,1,1,1,1,1,1,1,1,1,1,12,12,12,12,5,5,6,6,6,6,2,2,6,6,4,6,6,6,2,2,3,0,6,6,4,4,7,7,14,14,14,14,9,9,9,9,9,9,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,10,10,11,11,12,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,12,5,5,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,6,7,7,14,14,14,14,14,14,14,14,9,9,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,10,10,11,11,11,12,1,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,12,12,12,5,5,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,7,7,14,14,14,14,14,14,14,14,9,9,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,15,15,10,10,10,12,11,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,1,12,1,12,12,12,12,11,11,11,11,11,11,11,11,11,11,3,3,6,6,2,2,6,6,6,4,4,4,7,7,14,14,14,14,14,14,14,14,9,9,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,10,10,12,11,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,12,1,12,12,12,12,12,11,11,11,11,11,11,11,11,11,11,3,13,6,6,2,2,6,6,4,6,4,4,7,7,14,14,14,14,14,14,14,14,9,9,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,15,10,10,11,11,12,12,1,1,1,1,1,1,1,1,1,1,1,1,12,1,12,1,12,12,5,5,5,5,5,5,5,5,5,5,5,5,2,5,2,2,2,2,2,2,2,2,2,2,2,2,7,7,14,14,14,14,14,14,9,9,9,9,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,10,10,10,11,11,12,12,12,12,1,1,1,1,1,1,1,1,1,1,1,12,1,1,12,12,5,5,5,5,5,5,5,5,5,5,5,5,5,2,2,2,2,2,2,2,2,2,2,2,2,2,7,7,14,14,14,14,14,14,9,9,9,9,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,15,10,10,12,11,12,1,1,1,1,1,1,1,1,1,1,1,1,1,12,1,6,6,6,6,5,5,0,0,0,0,0,0,0,0,0,0,0,8,0,0,0,0,0,0,0,0,3,3,3,3,3,6,7,7,14,14,14,14,9,9,14,14,9,9,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,15,10,10,12,11,1,12,1,1,1,1,1,1,1,1,1,1,1,1,1,12,6,6,6,6,5,5,3,0,0,0,0,8,0,0,0,8,0,8,0,0,0,0,3,0,3,8,0,0,3,3,3,3,7,7,14,14,14,14,9,9,14,14,9,9,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,10,10,11,11,12,12,12,1,1,1,1,1,1,1,1,1,1,1,12,1,12,1,6,6,8,0,2,2,0,3,6,6,6,6,8,0,6,6,6,6,8,8,8,8,6,6,6,6,0,0,6,6,4,4,7,7,14,14,9,9,14,14,9,9,9,9,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,10,15,11,11,11,12,1,12,1,1,1,1,1,1,1,1,1,1,1,12,1,12,6,3,3,0,2,2,3,0,6,6,6,6,8,0,6,6,6,6,8,8,8,8,6,6,6,6,8,0,6,6,4,6,7,7,14,14,9,9,14,14,9,9,9,9,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,10,10,11,11,12,12,1,1,1,1,1,1,1,1,1,1,1,1,12,1,12,12,6,6,0,3,5,2,0,0,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,0,3,3,3,7,7,9,9,9,9,14,14,14,14,9,9,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,10,10,11,11,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,12,12,12,6,6,0,0,2,5,0,0,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,3,0,3,6,9,7,9,9,9,9,14,14,14,14,9,9,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,10,10,10,12,11,12,1,1,1,1,1,1,1,1,1,1,1,1,1,12,1,12,12,5,5,5,5,5,2,0,0,6,6,6,6,8,8,6,6,6,6,8,8,8,8,6,6,6,6,8,8,6,6,6,6,3,3,7,7,9,7,9,9,14,14,14,14,9,9,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,10,10,11,11,1,12,1,1,1,1,1,1,1,1,1,1,1,1,1,12,12,12,5,5,5,5,2,5,0,0,6,6,6,6,8,8,6,6,6,6,8,8,8,8,6,3,6,6,8,8,6,6,6,6,3,3,7,7,9,9,9,9,14,14,14,14,9,9,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,10,10,11,11,12,1,1,1,1,1,1,1,1,1,1,1,1,1,12,1,12,12,5,5,0,3,0,0,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,3,3,3,6,9,7,14,14,14,14,14,14,14,14,9,9,14,14,14),
(15,15,15,15,15,15,15,15,15,15,10,10,10,11,11,1,12,1,1,1,1,1,1,1,1,1,1,1,1,1,12,12,12,5,5,3,0,0,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,3,3,3,3,9,7,14,14,14,14,14,14,14,14,9,9,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,10,10,11,11,12,12,1,1,1,1,1,1,1,1,1,1,1,1,12,1,12,12,5,5,0,0,6,6,0,0,6,6,6,6,8,0,6,6,6,6,8,8,8,8,6,6,6,6,8,0,6,6,6,6,3,3,4,4,9,7,14,14,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,10,10,11,11,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,12,12,12,5,5,3,3,6,6,0,0,6,6,6,6,8,0,6,6,6,6,8,8,8,8,6,6,6,6,8,0,6,6,6,6,0,3,4,4,7,7,14,14,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,10,10,11,11,11,12,12,1,1,1,1,1,1,1,1,1,1,1,12,1,12,12,5,5,0,0,0,3,0,0,0,3,8,3,0,3,0,3,8,3,8,0,0,0,0,3,8,3,0,3,0,3,0,3,3,3,7,7,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,10,15,11,12,12,12,1,12,1,1,1,1,1,1,1,1,1,1,1,12,12,12,5,5,8,0,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,3,3,6,7,7,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,15,10,10,12,11,12,1,1,1,1,1,1,1,1,1,1,1,12,1,12,12,5,5,5,5,5,5,5,5,2,2,2,2,2,2,2,2,2,2,5,2,5,2,5,2,2,2,2,2,2,2,2,2,2,2,9,7,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,10,10,10,12,11,1,12,1,1,1,1,1,1,1,1,1,1,1,12,12,12,5,5,5,5,5,5,5,5,2,2,2,2,2,2,2,2,2,2,2,5,2,5,2,5,2,2,2,2,2,2,2,2,2,2,9,9,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,15,10,10,11,11,11,12,12,1,1,1,1,1,1,1,1,1,1,1,12,1,12,1,12,12,12,12,11,12,2,2,6,6,2,2,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,4,4,4,4,9,7,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,15,10,10,11,12,12,12,1,12,1,1,1,1,1,1,1,1,1,1,1,12,12,12,12,12,12,12,12,11,2,2,6,6,2,2,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,4,4,4,4,9,7,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,10,10,12,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,12,1,12,1,12,12,12,12,5,5,3,3,2,2,3,0,3,3,0,0,0,0,0,0,0,0,0,0,3,3,3,6,7,7,7,9,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,15,15,10,10,10,1,11,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,12,1,12,12,12,12,12,5,2,0,3,2,2,0,3,0,0,8,8,0,8,0,0,0,8,0,8,3,3,3,3,7,7,9,9,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,10,10,12,11,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,1,12,12,5,5,5,2,2,5,3,0,0,0,6,6,6,6,8,8,6,6,6,6,3,3,3,6,7,7,14,14,9,9,14,14,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,10,2,11,12,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,12,12,5,5,5,5,5,2,0,0,0,0,6,6,6,6,8,8,6,6,6,6,3,3,3,3,7,7,14,14,9,9,14,14,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,15,15,10,10,10,12,11,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,1,12,12,11,12,5,5,0,0,8,8,8,8,8,8,8,8,8,8,8,0,3,3,7,7,14,14,14,14,9,9,14,14,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,15,15,10,10,10,1,11,1,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,12,12,12,11,5,5,0,0,8,8,8,8,8,8,8,8,8,8,8,8,3,3,7,7,14,14,14,14,9,9,14,14,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,15,10,10,1,11,1,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,1,12,12,5,5,0,0,8,8,6,6,6,6,8,8,6,6,6,6,3,3,7,7,14,14,14,14,14,14,9,9,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,15,10,10,11,11,12,12,1,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,12,12,5,5,8,0,8,8,6,3,6,6,8,8,6,6,6,6,3,3,7,7,14,14,14,14,14,14,9,9,14,14,14,14,14,14,14,14,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,10,15,11,11,11,12,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,1,12,12,5,5,8,8,8,8,8,8,8,8,8,8,8,8,8,0,3,3,7,7,14,14,14,14,14,14,9,9,14,14,14,14,14,14,9,9,14,14,14),
(15,15,15,15,15,15,15,15,15,15,15,15,10,11,11,11,11,1,12,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,12,12,12,5,5,8,8,8,8,8,8,8,8,8,8,8,8,8,0,3,3,7,7,14,14,14,14,14,14,9,9,14,14,14,14,14,14,9,9,14,14,14)
);


end package sprites;